
  // Send an 'all' synchronized to all PE's 
  // pe__sys__thisSyncnronized basically means all the streams in a PE are complete
  // The PE controller will move to a 'final' state once it receives sys__pe__allSynchronized
  assign  GenStackBus[0].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[1].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[2].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[3].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[4].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[5].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[6].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[7].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[8].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[9].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[10].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[11].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[12].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[13].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[14].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[15].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[16].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[17].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[18].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[19].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[20].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[21].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[22].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[23].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[24].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[25].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[26].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[27].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[28].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[29].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[30].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[31].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[32].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[33].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[34].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[35].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[36].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[37].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[38].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[39].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[40].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[41].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[42].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[43].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[44].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[45].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[46].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[47].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[48].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[49].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[50].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[51].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[52].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[53].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[54].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[55].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[56].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[57].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[58].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[59].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[60].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[61].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[62].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 

  assign  GenStackBus[63].sys__pe__allSynchronized = GenStackBus[0].pe__sys__thisSynchronized & 
                                   GenStackBus[1].pe__sys__thisSynchronized & 
                                   GenStackBus[2].pe__sys__thisSynchronized & 
                                   GenStackBus[3].pe__sys__thisSynchronized & 
                                   GenStackBus[4].pe__sys__thisSynchronized & 
                                   GenStackBus[5].pe__sys__thisSynchronized & 
                                   GenStackBus[6].pe__sys__thisSynchronized & 
                                   GenStackBus[7].pe__sys__thisSynchronized & 
                                   GenStackBus[8].pe__sys__thisSynchronized & 
                                   GenStackBus[9].pe__sys__thisSynchronized & 
                                   GenStackBus[10].pe__sys__thisSynchronized & 
                                   GenStackBus[11].pe__sys__thisSynchronized & 
                                   GenStackBus[12].pe__sys__thisSynchronized & 
                                   GenStackBus[13].pe__sys__thisSynchronized & 
                                   GenStackBus[14].pe__sys__thisSynchronized & 
                                   GenStackBus[15].pe__sys__thisSynchronized & 
                                   GenStackBus[16].pe__sys__thisSynchronized & 
                                   GenStackBus[17].pe__sys__thisSynchronized & 
                                   GenStackBus[18].pe__sys__thisSynchronized & 
                                   GenStackBus[19].pe__sys__thisSynchronized & 
                                   GenStackBus[20].pe__sys__thisSynchronized & 
                                   GenStackBus[21].pe__sys__thisSynchronized & 
                                   GenStackBus[22].pe__sys__thisSynchronized & 
                                   GenStackBus[23].pe__sys__thisSynchronized & 
                                   GenStackBus[24].pe__sys__thisSynchronized & 
                                   GenStackBus[25].pe__sys__thisSynchronized & 
                                   GenStackBus[26].pe__sys__thisSynchronized & 
                                   GenStackBus[27].pe__sys__thisSynchronized & 
                                   GenStackBus[28].pe__sys__thisSynchronized & 
                                   GenStackBus[29].pe__sys__thisSynchronized & 
                                   GenStackBus[30].pe__sys__thisSynchronized & 
                                   GenStackBus[31].pe__sys__thisSynchronized & 
                                   GenStackBus[32].pe__sys__thisSynchronized & 
                                   GenStackBus[33].pe__sys__thisSynchronized & 
                                   GenStackBus[34].pe__sys__thisSynchronized & 
                                   GenStackBus[35].pe__sys__thisSynchronized & 
                                   GenStackBus[36].pe__sys__thisSynchronized & 
                                   GenStackBus[37].pe__sys__thisSynchronized & 
                                   GenStackBus[38].pe__sys__thisSynchronized & 
                                   GenStackBus[39].pe__sys__thisSynchronized & 
                                   GenStackBus[40].pe__sys__thisSynchronized & 
                                   GenStackBus[41].pe__sys__thisSynchronized & 
                                   GenStackBus[42].pe__sys__thisSynchronized & 
                                   GenStackBus[43].pe__sys__thisSynchronized & 
                                   GenStackBus[44].pe__sys__thisSynchronized & 
                                   GenStackBus[45].pe__sys__thisSynchronized & 
                                   GenStackBus[46].pe__sys__thisSynchronized & 
                                   GenStackBus[47].pe__sys__thisSynchronized & 
                                   GenStackBus[48].pe__sys__thisSynchronized & 
                                   GenStackBus[49].pe__sys__thisSynchronized & 
                                   GenStackBus[50].pe__sys__thisSynchronized & 
                                   GenStackBus[51].pe__sys__thisSynchronized & 
                                   GenStackBus[52].pe__sys__thisSynchronized & 
                                   GenStackBus[53].pe__sys__thisSynchronized & 
                                   GenStackBus[54].pe__sys__thisSynchronized & 
                                   GenStackBus[55].pe__sys__thisSynchronized & 
                                   GenStackBus[56].pe__sys__thisSynchronized & 
                                   GenStackBus[57].pe__sys__thisSynchronized & 
                                   GenStackBus[58].pe__sys__thisSynchronized & 
                                   GenStackBus[59].pe__sys__thisSynchronized & 
                                   GenStackBus[60].pe__sys__thisSynchronized & 
                                   GenStackBus[61].pe__sys__thisSynchronized & 
                                   GenStackBus[62].pe__sys__thisSynchronized & 
                                   GenStackBus[63].pe__sys__thisSynchronized ; 
