
  // General control and status                                       
  assign    sys__pe0__allSynchronized     =    mgr0__sys__allSynchronized   ;
  assign    sys__mgr0__thisSynchronized   =    pe0__sys__thisSynchronized   ;
  assign    sys__mgr0__ready              =    pe0__sys__ready              ;
  assign    sys__mgr0__complete           =    pe0__sys__complete           ;

  // General control and status                                       
  assign    sys__pe1__allSynchronized     =    mgr1__sys__allSynchronized   ;
  assign    sys__mgr1__thisSynchronized   =    pe1__sys__thisSynchronized   ;
  assign    sys__mgr1__ready              =    pe1__sys__ready              ;
  assign    sys__mgr1__complete           =    pe1__sys__complete           ;

  // General control and status                                       
  assign    sys__pe2__allSynchronized     =    mgr2__sys__allSynchronized   ;
  assign    sys__mgr2__thisSynchronized   =    pe2__sys__thisSynchronized   ;
  assign    sys__mgr2__ready              =    pe2__sys__ready              ;
  assign    sys__mgr2__complete           =    pe2__sys__complete           ;

  // General control and status                                       
  assign    sys__pe3__allSynchronized     =    mgr3__sys__allSynchronized   ;
  assign    sys__mgr3__thisSynchronized   =    pe3__sys__thisSynchronized   ;
  assign    sys__mgr3__ready              =    pe3__sys__ready              ;
  assign    sys__mgr3__complete           =    pe3__sys__complete           ;
