
               // General control and status                                                 
               .sys__pe__peId                      ( sys__pe__peId                   ),      
               .sys__pe__allSynchronized           ( sys__pe__allSynchronized        ),      
               .pe__sys__thisSynchronized          ( pe__sys__thisSynchronized       ),      
               .pe__sys__ready                     ( pe__sys__ready                  ),      
               .pe__sys__complete                  ( pe__sys__complete               ),      