
            begin
                @vSysLane2PeArray[0][0].cb_test                                      ;
                vSysLane2PeArray [0][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][1].cb_test                                      ;
                vSysLane2PeArray [0][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][2].cb_test                                      ;
                vSysLane2PeArray [0][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][3].cb_test                                      ;
                vSysLane2PeArray [0][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][4].cb_test                                      ;
                vSysLane2PeArray [0][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][5].cb_test                                      ;
                vSysLane2PeArray [0][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][6].cb_test                                      ;
                vSysLane2PeArray [0][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][7].cb_test                                      ;
                vSysLane2PeArray [0][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][8].cb_test                                      ;
                vSysLane2PeArray [0][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][9].cb_test                                      ;
                vSysLane2PeArray [0][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][10].cb_test                                      ;
                vSysLane2PeArray [0][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][11].cb_test                                      ;
                vSysLane2PeArray [0][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][12].cb_test                                      ;
                vSysLane2PeArray [0][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][13].cb_test                                      ;
                vSysLane2PeArray [0][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][14].cb_test                                      ;
                vSysLane2PeArray [0][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][15].cb_test                                      ;
                vSysLane2PeArray [0][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][16].cb_test                                      ;
                vSysLane2PeArray [0][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][17].cb_test                                      ;
                vSysLane2PeArray [0][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][18].cb_test                                      ;
                vSysLane2PeArray [0][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][19].cb_test                                      ;
                vSysLane2PeArray [0][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][20].cb_test                                      ;
                vSysLane2PeArray [0][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][21].cb_test                                      ;
                vSysLane2PeArray [0][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][22].cb_test                                      ;
                vSysLane2PeArray [0][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][23].cb_test                                      ;
                vSysLane2PeArray [0][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][24].cb_test                                      ;
                vSysLane2PeArray [0][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][25].cb_test                                      ;
                vSysLane2PeArray [0][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][26].cb_test                                      ;
                vSysLane2PeArray [0][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][27].cb_test                                      ;
                vSysLane2PeArray [0][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][28].cb_test                                      ;
                vSysLane2PeArray [0][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][29].cb_test                                      ;
                vSysLane2PeArray [0][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][30].cb_test                                      ;
                vSysLane2PeArray [0][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[0][31].cb_test                                      ;
                vSysLane2PeArray [0][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [0][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSysLane2PeArray[1][0].cb_test                                      ;
                vSysLane2PeArray [1][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][1].cb_test                                      ;
                vSysLane2PeArray [1][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][2].cb_test                                      ;
                vSysLane2PeArray [1][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][3].cb_test                                      ;
                vSysLane2PeArray [1][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][4].cb_test                                      ;
                vSysLane2PeArray [1][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][5].cb_test                                      ;
                vSysLane2PeArray [1][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][6].cb_test                                      ;
                vSysLane2PeArray [1][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][7].cb_test                                      ;
                vSysLane2PeArray [1][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][8].cb_test                                      ;
                vSysLane2PeArray [1][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][9].cb_test                                      ;
                vSysLane2PeArray [1][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][10].cb_test                                      ;
                vSysLane2PeArray [1][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][11].cb_test                                      ;
                vSysLane2PeArray [1][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][12].cb_test                                      ;
                vSysLane2PeArray [1][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][13].cb_test                                      ;
                vSysLane2PeArray [1][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][14].cb_test                                      ;
                vSysLane2PeArray [1][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][15].cb_test                                      ;
                vSysLane2PeArray [1][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][16].cb_test                                      ;
                vSysLane2PeArray [1][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][17].cb_test                                      ;
                vSysLane2PeArray [1][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][18].cb_test                                      ;
                vSysLane2PeArray [1][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][19].cb_test                                      ;
                vSysLane2PeArray [1][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][20].cb_test                                      ;
                vSysLane2PeArray [1][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][21].cb_test                                      ;
                vSysLane2PeArray [1][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][22].cb_test                                      ;
                vSysLane2PeArray [1][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][23].cb_test                                      ;
                vSysLane2PeArray [1][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][24].cb_test                                      ;
                vSysLane2PeArray [1][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][25].cb_test                                      ;
                vSysLane2PeArray [1][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][26].cb_test                                      ;
                vSysLane2PeArray [1][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][27].cb_test                                      ;
                vSysLane2PeArray [1][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][28].cb_test                                      ;
                vSysLane2PeArray [1][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][29].cb_test                                      ;
                vSysLane2PeArray [1][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][30].cb_test                                      ;
                vSysLane2PeArray [1][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[1][31].cb_test                                      ;
                vSysLane2PeArray [1][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [1][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSysLane2PeArray[2][0].cb_test                                      ;
                vSysLane2PeArray [2][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][1].cb_test                                      ;
                vSysLane2PeArray [2][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][2].cb_test                                      ;
                vSysLane2PeArray [2][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][3].cb_test                                      ;
                vSysLane2PeArray [2][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][4].cb_test                                      ;
                vSysLane2PeArray [2][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][5].cb_test                                      ;
                vSysLane2PeArray [2][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][6].cb_test                                      ;
                vSysLane2PeArray [2][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][7].cb_test                                      ;
                vSysLane2PeArray [2][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][8].cb_test                                      ;
                vSysLane2PeArray [2][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][9].cb_test                                      ;
                vSysLane2PeArray [2][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][10].cb_test                                      ;
                vSysLane2PeArray [2][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][11].cb_test                                      ;
                vSysLane2PeArray [2][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][12].cb_test                                      ;
                vSysLane2PeArray [2][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][13].cb_test                                      ;
                vSysLane2PeArray [2][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][14].cb_test                                      ;
                vSysLane2PeArray [2][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][15].cb_test                                      ;
                vSysLane2PeArray [2][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][16].cb_test                                      ;
                vSysLane2PeArray [2][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][17].cb_test                                      ;
                vSysLane2PeArray [2][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][18].cb_test                                      ;
                vSysLane2PeArray [2][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][19].cb_test                                      ;
                vSysLane2PeArray [2][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][20].cb_test                                      ;
                vSysLane2PeArray [2][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][21].cb_test                                      ;
                vSysLane2PeArray [2][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][22].cb_test                                      ;
                vSysLane2PeArray [2][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][23].cb_test                                      ;
                vSysLane2PeArray [2][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][24].cb_test                                      ;
                vSysLane2PeArray [2][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][25].cb_test                                      ;
                vSysLane2PeArray [2][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][26].cb_test                                      ;
                vSysLane2PeArray [2][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][27].cb_test                                      ;
                vSysLane2PeArray [2][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][28].cb_test                                      ;
                vSysLane2PeArray [2][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][29].cb_test                                      ;
                vSysLane2PeArray [2][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][30].cb_test                                      ;
                vSysLane2PeArray [2][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[2][31].cb_test                                      ;
                vSysLane2PeArray [2][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [2][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSysLane2PeArray[3][0].cb_test                                      ;
                vSysLane2PeArray [3][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][1].cb_test                                      ;
                vSysLane2PeArray [3][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][2].cb_test                                      ;
                vSysLane2PeArray [3][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][3].cb_test                                      ;
                vSysLane2PeArray [3][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][4].cb_test                                      ;
                vSysLane2PeArray [3][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][5].cb_test                                      ;
                vSysLane2PeArray [3][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][6].cb_test                                      ;
                vSysLane2PeArray [3][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][7].cb_test                                      ;
                vSysLane2PeArray [3][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][8].cb_test                                      ;
                vSysLane2PeArray [3][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][9].cb_test                                      ;
                vSysLane2PeArray [3][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][10].cb_test                                      ;
                vSysLane2PeArray [3][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][11].cb_test                                      ;
                vSysLane2PeArray [3][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][12].cb_test                                      ;
                vSysLane2PeArray [3][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][13].cb_test                                      ;
                vSysLane2PeArray [3][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][14].cb_test                                      ;
                vSysLane2PeArray [3][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][15].cb_test                                      ;
                vSysLane2PeArray [3][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][16].cb_test                                      ;
                vSysLane2PeArray [3][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][17].cb_test                                      ;
                vSysLane2PeArray [3][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][18].cb_test                                      ;
                vSysLane2PeArray [3][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][19].cb_test                                      ;
                vSysLane2PeArray [3][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][20].cb_test                                      ;
                vSysLane2PeArray [3][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][21].cb_test                                      ;
                vSysLane2PeArray [3][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][22].cb_test                                      ;
                vSysLane2PeArray [3][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][23].cb_test                                      ;
                vSysLane2PeArray [3][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][24].cb_test                                      ;
                vSysLane2PeArray [3][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][25].cb_test                                      ;
                vSysLane2PeArray [3][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][26].cb_test                                      ;
                vSysLane2PeArray [3][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][27].cb_test                                      ;
                vSysLane2PeArray [3][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][28].cb_test                                      ;
                vSysLane2PeArray [3][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][29].cb_test                                      ;
                vSysLane2PeArray [3][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][30].cb_test                                      ;
                vSysLane2PeArray [3][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSysLane2PeArray[3][31].cb_test                                      ;
                vSysLane2PeArray [3][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSysLane2PeArray [3][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
