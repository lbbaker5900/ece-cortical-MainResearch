
    wire                                           stu__mgr0__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr0__cntl           ;
    wire                                           mgr0__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr0__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr0__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr0__oob_data       ;

    wire                                           stu__mgr1__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr1__cntl           ;
    wire                                           mgr1__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr1__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr1__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr1__oob_data       ;

    wire                                           stu__mgr2__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr2__cntl           ;
    wire                                           mgr2__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr2__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr2__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr2__oob_data       ;

    wire                                           stu__mgr3__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr3__cntl           ;
    wire                                           mgr3__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr3__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr3__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr3__oob_data       ;

    wire                                           stu__mgr4__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr4__cntl           ;
    wire                                           mgr4__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr4__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr4__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr4__oob_data       ;

    wire                                           stu__mgr5__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr5__cntl           ;
    wire                                           mgr5__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr5__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr5__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr5__oob_data       ;

    wire                                           stu__mgr6__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr6__cntl           ;
    wire                                           mgr6__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr6__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr6__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr6__oob_data       ;

    wire                                           stu__mgr7__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr7__cntl           ;
    wire                                           mgr7__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr7__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr7__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr7__oob_data       ;

    wire                                           stu__mgr8__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr8__cntl           ;
    wire                                           mgr8__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr8__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr8__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr8__oob_data       ;

    wire                                           stu__mgr9__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr9__cntl           ;
    wire                                           mgr9__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr9__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr9__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr9__oob_data       ;

    wire                                           stu__mgr10__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr10__cntl           ;
    wire                                           mgr10__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr10__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr10__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr10__oob_data       ;

    wire                                           stu__mgr11__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr11__cntl           ;
    wire                                           mgr11__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr11__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr11__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr11__oob_data       ;

    wire                                           stu__mgr12__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr12__cntl           ;
    wire                                           mgr12__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr12__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr12__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr12__oob_data       ;

    wire                                           stu__mgr13__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr13__cntl           ;
    wire                                           mgr13__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr13__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr13__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr13__oob_data       ;

    wire                                           stu__mgr14__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr14__cntl           ;
    wire                                           mgr14__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr14__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr14__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr14__oob_data       ;

    wire                                           stu__mgr15__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr15__cntl           ;
    wire                                           mgr15__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr15__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr15__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr15__oob_data       ;

    wire                                           stu__mgr16__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr16__cntl           ;
    wire                                           mgr16__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr16__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr16__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr16__oob_data       ;

    wire                                           stu__mgr17__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr17__cntl           ;
    wire                                           mgr17__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr17__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr17__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr17__oob_data       ;

    wire                                           stu__mgr18__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr18__cntl           ;
    wire                                           mgr18__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr18__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr18__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr18__oob_data       ;

    wire                                           stu__mgr19__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr19__cntl           ;
    wire                                           mgr19__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr19__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr19__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr19__oob_data       ;

    wire                                           stu__mgr20__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr20__cntl           ;
    wire                                           mgr20__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr20__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr20__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr20__oob_data       ;

    wire                                           stu__mgr21__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr21__cntl           ;
    wire                                           mgr21__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr21__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr21__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr21__oob_data       ;

    wire                                           stu__mgr22__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr22__cntl           ;
    wire                                           mgr22__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr22__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr22__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr22__oob_data       ;

    wire                                           stu__mgr23__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr23__cntl           ;
    wire                                           mgr23__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr23__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr23__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr23__oob_data       ;

    wire                                           stu__mgr24__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr24__cntl           ;
    wire                                           mgr24__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr24__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr24__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr24__oob_data       ;

    wire                                           stu__mgr25__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr25__cntl           ;
    wire                                           mgr25__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr25__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr25__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr25__oob_data       ;

    wire                                           stu__mgr26__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr26__cntl           ;
    wire                                           mgr26__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr26__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr26__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr26__oob_data       ;

    wire                                           stu__mgr27__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr27__cntl           ;
    wire                                           mgr27__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr27__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr27__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr27__oob_data       ;

    wire                                           stu__mgr28__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr28__cntl           ;
    wire                                           mgr28__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr28__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr28__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr28__oob_data       ;

    wire                                           stu__mgr29__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr29__cntl           ;
    wire                                           mgr29__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr29__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr29__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr29__oob_data       ;

    wire                                           stu__mgr30__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr30__cntl           ;
    wire                                           mgr30__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr30__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr30__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr30__oob_data       ;

    wire                                           stu__mgr31__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr31__cntl           ;
    wire                                           mgr31__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr31__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr31__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr31__oob_data       ;

    wire                                           stu__mgr32__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr32__cntl           ;
    wire                                           mgr32__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr32__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr32__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr32__oob_data       ;

    wire                                           stu__mgr33__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr33__cntl           ;
    wire                                           mgr33__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr33__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr33__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr33__oob_data       ;

    wire                                           stu__mgr34__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr34__cntl           ;
    wire                                           mgr34__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr34__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr34__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr34__oob_data       ;

    wire                                           stu__mgr35__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr35__cntl           ;
    wire                                           mgr35__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr35__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr35__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr35__oob_data       ;

    wire                                           stu__mgr36__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr36__cntl           ;
    wire                                           mgr36__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr36__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr36__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr36__oob_data       ;

    wire                                           stu__mgr37__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr37__cntl           ;
    wire                                           mgr37__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr37__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr37__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr37__oob_data       ;

    wire                                           stu__mgr38__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr38__cntl           ;
    wire                                           mgr38__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr38__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr38__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr38__oob_data       ;

    wire                                           stu__mgr39__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr39__cntl           ;
    wire                                           mgr39__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr39__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr39__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr39__oob_data       ;

    wire                                           stu__mgr40__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr40__cntl           ;
    wire                                           mgr40__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr40__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr40__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr40__oob_data       ;

    wire                                           stu__mgr41__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr41__cntl           ;
    wire                                           mgr41__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr41__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr41__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr41__oob_data       ;

    wire                                           stu__mgr42__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr42__cntl           ;
    wire                                           mgr42__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr42__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr42__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr42__oob_data       ;

    wire                                           stu__mgr43__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr43__cntl           ;
    wire                                           mgr43__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr43__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr43__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr43__oob_data       ;

    wire                                           stu__mgr44__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr44__cntl           ;
    wire                                           mgr44__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr44__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr44__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr44__oob_data       ;

    wire                                           stu__mgr45__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr45__cntl           ;
    wire                                           mgr45__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr45__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr45__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr45__oob_data       ;

    wire                                           stu__mgr46__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr46__cntl           ;
    wire                                           mgr46__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr46__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr46__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr46__oob_data       ;

    wire                                           stu__mgr47__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr47__cntl           ;
    wire                                           mgr47__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr47__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr47__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr47__oob_data       ;

    wire                                           stu__mgr48__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr48__cntl           ;
    wire                                           mgr48__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr48__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr48__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr48__oob_data       ;

    wire                                           stu__mgr49__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr49__cntl           ;
    wire                                           mgr49__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr49__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr49__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr49__oob_data       ;

    wire                                           stu__mgr50__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr50__cntl           ;
    wire                                           mgr50__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr50__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr50__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr50__oob_data       ;

    wire                                           stu__mgr51__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr51__cntl           ;
    wire                                           mgr51__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr51__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr51__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr51__oob_data       ;

    wire                                           stu__mgr52__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr52__cntl           ;
    wire                                           mgr52__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr52__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr52__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr52__oob_data       ;

    wire                                           stu__mgr53__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr53__cntl           ;
    wire                                           mgr53__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr53__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr53__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr53__oob_data       ;

    wire                                           stu__mgr54__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr54__cntl           ;
    wire                                           mgr54__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr54__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr54__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr54__oob_data       ;

    wire                                           stu__mgr55__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr55__cntl           ;
    wire                                           mgr55__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr55__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr55__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr55__oob_data       ;

    wire                                           stu__mgr56__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr56__cntl           ;
    wire                                           mgr56__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr56__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr56__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr56__oob_data       ;

    wire                                           stu__mgr57__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr57__cntl           ;
    wire                                           mgr57__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr57__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr57__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr57__oob_data       ;

    wire                                           stu__mgr58__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr58__cntl           ;
    wire                                           mgr58__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr58__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr58__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr58__oob_data       ;

    wire                                           stu__mgr59__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr59__cntl           ;
    wire                                           mgr59__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr59__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr59__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr59__oob_data       ;

    wire                                           stu__mgr60__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr60__cntl           ;
    wire                                           mgr60__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr60__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr60__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr60__oob_data       ;

    wire                                           stu__mgr61__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr61__cntl           ;
    wire                                           mgr61__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr61__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr61__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr61__oob_data       ;

    wire                                           stu__mgr62__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr62__cntl           ;
    wire                                           mgr62__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr62__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr62__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr62__oob_data       ;

    wire                                           stu__mgr63__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr63__cntl           ;
    wire                                           mgr63__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr63__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr63__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr63__oob_data       ;

