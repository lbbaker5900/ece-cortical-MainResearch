
  wire                                          dma__memc__lane0_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane0_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane0_write_data0            ;
  wire                                          memc__dma__lane0_write_ready0           ;
  wire                                          dma__memc__lane0_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane0_read_address0          ;
  wire                                          dma__memc__lane0_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane0_read_data0             ;
  wire                                          memc__dma__lane0_read_data_valid0       ;
  wire                                          memc__dma__lane0_read_ready0            ;
  wire                                          dma__memc__lane1_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane1_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane1_write_data0            ;
  wire                                          memc__dma__lane1_write_ready0           ;
  wire                                          dma__memc__lane1_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane1_read_address0          ;
  wire                                          dma__memc__lane1_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane1_read_data0             ;
  wire                                          memc__dma__lane1_read_data_valid0       ;
  wire                                          memc__dma__lane1_read_ready0            ;
  wire                                          dma__memc__lane2_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane2_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane2_write_data0            ;
  wire                                          memc__dma__lane2_write_ready0           ;
  wire                                          dma__memc__lane2_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane2_read_address0          ;
  wire                                          dma__memc__lane2_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane2_read_data0             ;
  wire                                          memc__dma__lane2_read_data_valid0       ;
  wire                                          memc__dma__lane2_read_ready0            ;
  wire                                          dma__memc__lane3_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane3_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane3_write_data0            ;
  wire                                          memc__dma__lane3_write_ready0           ;
  wire                                          dma__memc__lane3_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane3_read_address0          ;
  wire                                          dma__memc__lane3_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane3_read_data0             ;
  wire                                          memc__dma__lane3_read_data_valid0       ;
  wire                                          memc__dma__lane3_read_ready0            ;
  wire                                          dma__memc__lane4_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane4_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane4_write_data0            ;
  wire                                          memc__dma__lane4_write_ready0           ;
  wire                                          dma__memc__lane4_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane4_read_address0          ;
  wire                                          dma__memc__lane4_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane4_read_data0             ;
  wire                                          memc__dma__lane4_read_data_valid0       ;
  wire                                          memc__dma__lane4_read_ready0            ;
  wire                                          dma__memc__lane5_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane5_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane5_write_data0            ;
  wire                                          memc__dma__lane5_write_ready0           ;
  wire                                          dma__memc__lane5_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane5_read_address0          ;
  wire                                          dma__memc__lane5_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane5_read_data0             ;
  wire                                          memc__dma__lane5_read_data_valid0       ;
  wire                                          memc__dma__lane5_read_ready0            ;
  wire                                          dma__memc__lane6_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane6_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane6_write_data0            ;
  wire                                          memc__dma__lane6_write_ready0           ;
  wire                                          dma__memc__lane6_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane6_read_address0          ;
  wire                                          dma__memc__lane6_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane6_read_data0             ;
  wire                                          memc__dma__lane6_read_data_valid0       ;
  wire                                          memc__dma__lane6_read_ready0            ;
  wire                                          dma__memc__lane7_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane7_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane7_write_data0            ;
  wire                                          memc__dma__lane7_write_ready0           ;
  wire                                          dma__memc__lane7_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane7_read_address0          ;
  wire                                          dma__memc__lane7_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane7_read_data0             ;
  wire                                          memc__dma__lane7_read_data_valid0       ;
  wire                                          memc__dma__lane7_read_ready0            ;
  wire                                          dma__memc__lane8_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane8_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane8_write_data0            ;
  wire                                          memc__dma__lane8_write_ready0           ;
  wire                                          dma__memc__lane8_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane8_read_address0          ;
  wire                                          dma__memc__lane8_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane8_read_data0             ;
  wire                                          memc__dma__lane8_read_data_valid0       ;
  wire                                          memc__dma__lane8_read_ready0            ;
  wire                                          dma__memc__lane9_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane9_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane9_write_data0            ;
  wire                                          memc__dma__lane9_write_ready0           ;
  wire                                          dma__memc__lane9_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane9_read_address0          ;
  wire                                          dma__memc__lane9_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane9_read_data0             ;
  wire                                          memc__dma__lane9_read_data_valid0       ;
  wire                                          memc__dma__lane9_read_ready0            ;
  wire                                          dma__memc__lane10_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane10_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane10_write_data0            ;
  wire                                          memc__dma__lane10_write_ready0           ;
  wire                                          dma__memc__lane10_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane10_read_address0          ;
  wire                                          dma__memc__lane10_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane10_read_data0             ;
  wire                                          memc__dma__lane10_read_data_valid0       ;
  wire                                          memc__dma__lane10_read_ready0            ;
  wire                                          dma__memc__lane11_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane11_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane11_write_data0            ;
  wire                                          memc__dma__lane11_write_ready0           ;
  wire                                          dma__memc__lane11_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane11_read_address0          ;
  wire                                          dma__memc__lane11_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane11_read_data0             ;
  wire                                          memc__dma__lane11_read_data_valid0       ;
  wire                                          memc__dma__lane11_read_ready0            ;
  wire                                          dma__memc__lane12_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane12_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane12_write_data0            ;
  wire                                          memc__dma__lane12_write_ready0           ;
  wire                                          dma__memc__lane12_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane12_read_address0          ;
  wire                                          dma__memc__lane12_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane12_read_data0             ;
  wire                                          memc__dma__lane12_read_data_valid0       ;
  wire                                          memc__dma__lane12_read_ready0            ;
  wire                                          dma__memc__lane13_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane13_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane13_write_data0            ;
  wire                                          memc__dma__lane13_write_ready0           ;
  wire                                          dma__memc__lane13_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane13_read_address0          ;
  wire                                          dma__memc__lane13_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane13_read_data0             ;
  wire                                          memc__dma__lane13_read_data_valid0       ;
  wire                                          memc__dma__lane13_read_ready0            ;
  wire                                          dma__memc__lane14_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane14_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane14_write_data0            ;
  wire                                          memc__dma__lane14_write_ready0           ;
  wire                                          dma__memc__lane14_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane14_read_address0          ;
  wire                                          dma__memc__lane14_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane14_read_data0             ;
  wire                                          memc__dma__lane14_read_data_valid0       ;
  wire                                          memc__dma__lane14_read_ready0            ;
  wire                                          dma__memc__lane15_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane15_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane15_write_data0            ;
  wire                                          memc__dma__lane15_write_ready0           ;
  wire                                          dma__memc__lane15_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane15_read_address0          ;
  wire                                          dma__memc__lane15_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane15_read_data0             ;
  wire                                          memc__dma__lane15_read_data_valid0       ;
  wire                                          memc__dma__lane15_read_ready0            ;
  wire                                          dma__memc__lane16_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane16_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane16_write_data0            ;
  wire                                          memc__dma__lane16_write_ready0           ;
  wire                                          dma__memc__lane16_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane16_read_address0          ;
  wire                                          dma__memc__lane16_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane16_read_data0             ;
  wire                                          memc__dma__lane16_read_data_valid0       ;
  wire                                          memc__dma__lane16_read_ready0            ;
  wire                                          dma__memc__lane17_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane17_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane17_write_data0            ;
  wire                                          memc__dma__lane17_write_ready0           ;
  wire                                          dma__memc__lane17_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane17_read_address0          ;
  wire                                          dma__memc__lane17_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane17_read_data0             ;
  wire                                          memc__dma__lane17_read_data_valid0       ;
  wire                                          memc__dma__lane17_read_ready0            ;
  wire                                          dma__memc__lane18_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane18_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane18_write_data0            ;
  wire                                          memc__dma__lane18_write_ready0           ;
  wire                                          dma__memc__lane18_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane18_read_address0          ;
  wire                                          dma__memc__lane18_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane18_read_data0             ;
  wire                                          memc__dma__lane18_read_data_valid0       ;
  wire                                          memc__dma__lane18_read_ready0            ;
  wire                                          dma__memc__lane19_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane19_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane19_write_data0            ;
  wire                                          memc__dma__lane19_write_ready0           ;
  wire                                          dma__memc__lane19_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane19_read_address0          ;
  wire                                          dma__memc__lane19_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane19_read_data0             ;
  wire                                          memc__dma__lane19_read_data_valid0       ;
  wire                                          memc__dma__lane19_read_ready0            ;
  wire                                          dma__memc__lane20_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane20_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane20_write_data0            ;
  wire                                          memc__dma__lane20_write_ready0           ;
  wire                                          dma__memc__lane20_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane20_read_address0          ;
  wire                                          dma__memc__lane20_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane20_read_data0             ;
  wire                                          memc__dma__lane20_read_data_valid0       ;
  wire                                          memc__dma__lane20_read_ready0            ;
  wire                                          dma__memc__lane21_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane21_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane21_write_data0            ;
  wire                                          memc__dma__lane21_write_ready0           ;
  wire                                          dma__memc__lane21_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane21_read_address0          ;
  wire                                          dma__memc__lane21_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane21_read_data0             ;
  wire                                          memc__dma__lane21_read_data_valid0       ;
  wire                                          memc__dma__lane21_read_ready0            ;
  wire                                          dma__memc__lane22_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane22_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane22_write_data0            ;
  wire                                          memc__dma__lane22_write_ready0           ;
  wire                                          dma__memc__lane22_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane22_read_address0          ;
  wire                                          dma__memc__lane22_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane22_read_data0             ;
  wire                                          memc__dma__lane22_read_data_valid0       ;
  wire                                          memc__dma__lane22_read_ready0            ;
  wire                                          dma__memc__lane23_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane23_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane23_write_data0            ;
  wire                                          memc__dma__lane23_write_ready0           ;
  wire                                          dma__memc__lane23_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane23_read_address0          ;
  wire                                          dma__memc__lane23_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane23_read_data0             ;
  wire                                          memc__dma__lane23_read_data_valid0       ;
  wire                                          memc__dma__lane23_read_ready0            ;
  wire                                          dma__memc__lane24_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane24_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane24_write_data0            ;
  wire                                          memc__dma__lane24_write_ready0           ;
  wire                                          dma__memc__lane24_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane24_read_address0          ;
  wire                                          dma__memc__lane24_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane24_read_data0             ;
  wire                                          memc__dma__lane24_read_data_valid0       ;
  wire                                          memc__dma__lane24_read_ready0            ;
  wire                                          dma__memc__lane25_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane25_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane25_write_data0            ;
  wire                                          memc__dma__lane25_write_ready0           ;
  wire                                          dma__memc__lane25_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane25_read_address0          ;
  wire                                          dma__memc__lane25_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane25_read_data0             ;
  wire                                          memc__dma__lane25_read_data_valid0       ;
  wire                                          memc__dma__lane25_read_ready0            ;
  wire                                          dma__memc__lane26_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane26_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane26_write_data0            ;
  wire                                          memc__dma__lane26_write_ready0           ;
  wire                                          dma__memc__lane26_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane26_read_address0          ;
  wire                                          dma__memc__lane26_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane26_read_data0             ;
  wire                                          memc__dma__lane26_read_data_valid0       ;
  wire                                          memc__dma__lane26_read_ready0            ;
  wire                                          dma__memc__lane27_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane27_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane27_write_data0            ;
  wire                                          memc__dma__lane27_write_ready0           ;
  wire                                          dma__memc__lane27_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane27_read_address0          ;
  wire                                          dma__memc__lane27_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane27_read_data0             ;
  wire                                          memc__dma__lane27_read_data_valid0       ;
  wire                                          memc__dma__lane27_read_ready0            ;
  wire                                          dma__memc__lane28_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane28_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane28_write_data0            ;
  wire                                          memc__dma__lane28_write_ready0           ;
  wire                                          dma__memc__lane28_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane28_read_address0          ;
  wire                                          dma__memc__lane28_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane28_read_data0             ;
  wire                                          memc__dma__lane28_read_data_valid0       ;
  wire                                          memc__dma__lane28_read_ready0            ;
  wire                                          dma__memc__lane29_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane29_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane29_write_data0            ;
  wire                                          memc__dma__lane29_write_ready0           ;
  wire                                          dma__memc__lane29_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane29_read_address0          ;
  wire                                          dma__memc__lane29_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane29_read_data0             ;
  wire                                          memc__dma__lane29_read_data_valid0       ;
  wire                                          memc__dma__lane29_read_ready0            ;
  wire                                          dma__memc__lane30_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane30_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane30_write_data0            ;
  wire                                          memc__dma__lane30_write_ready0           ;
  wire                                          dma__memc__lane30_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane30_read_address0          ;
  wire                                          dma__memc__lane30_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane30_read_data0             ;
  wire                                          memc__dma__lane30_read_data_valid0       ;
  wire                                          memc__dma__lane30_read_ready0            ;
  wire                                          dma__memc__lane31_write_valid0           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane31_write_address0         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane31_write_data0            ;
  wire                                          memc__dma__lane31_write_ready0           ;
  wire                                          dma__memc__lane31_read_valid0            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane31_read_address0          ;
  wire                                          dma__memc__lane31_read_pause0            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane31_read_data0             ;
  wire                                          memc__dma__lane31_read_data_valid0       ;
  wire                                          memc__dma__lane31_read_ready0            ;

  wire                                          dma__memc__lane0_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane0_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane0_write_data1            ;
  wire                                          memc__dma__lane0_write_ready1           ;
  wire                                          dma__memc__lane0_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane0_read_address1          ;
  wire                                          dma__memc__lane0_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane0_read_data1             ;
  wire                                          memc__dma__lane0_read_data_valid1       ;
  wire                                          memc__dma__lane0_read_ready1            ;
  wire                                          dma__memc__lane1_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane1_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane1_write_data1            ;
  wire                                          memc__dma__lane1_write_ready1           ;
  wire                                          dma__memc__lane1_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane1_read_address1          ;
  wire                                          dma__memc__lane1_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane1_read_data1             ;
  wire                                          memc__dma__lane1_read_data_valid1       ;
  wire                                          memc__dma__lane1_read_ready1            ;
  wire                                          dma__memc__lane2_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane2_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane2_write_data1            ;
  wire                                          memc__dma__lane2_write_ready1           ;
  wire                                          dma__memc__lane2_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane2_read_address1          ;
  wire                                          dma__memc__lane2_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane2_read_data1             ;
  wire                                          memc__dma__lane2_read_data_valid1       ;
  wire                                          memc__dma__lane2_read_ready1            ;
  wire                                          dma__memc__lane3_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane3_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane3_write_data1            ;
  wire                                          memc__dma__lane3_write_ready1           ;
  wire                                          dma__memc__lane3_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane3_read_address1          ;
  wire                                          dma__memc__lane3_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane3_read_data1             ;
  wire                                          memc__dma__lane3_read_data_valid1       ;
  wire                                          memc__dma__lane3_read_ready1            ;
  wire                                          dma__memc__lane4_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane4_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane4_write_data1            ;
  wire                                          memc__dma__lane4_write_ready1           ;
  wire                                          dma__memc__lane4_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane4_read_address1          ;
  wire                                          dma__memc__lane4_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane4_read_data1             ;
  wire                                          memc__dma__lane4_read_data_valid1       ;
  wire                                          memc__dma__lane4_read_ready1            ;
  wire                                          dma__memc__lane5_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane5_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane5_write_data1            ;
  wire                                          memc__dma__lane5_write_ready1           ;
  wire                                          dma__memc__lane5_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane5_read_address1          ;
  wire                                          dma__memc__lane5_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane5_read_data1             ;
  wire                                          memc__dma__lane5_read_data_valid1       ;
  wire                                          memc__dma__lane5_read_ready1            ;
  wire                                          dma__memc__lane6_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane6_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane6_write_data1            ;
  wire                                          memc__dma__lane6_write_ready1           ;
  wire                                          dma__memc__lane6_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane6_read_address1          ;
  wire                                          dma__memc__lane6_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane6_read_data1             ;
  wire                                          memc__dma__lane6_read_data_valid1       ;
  wire                                          memc__dma__lane6_read_ready1            ;
  wire                                          dma__memc__lane7_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane7_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane7_write_data1            ;
  wire                                          memc__dma__lane7_write_ready1           ;
  wire                                          dma__memc__lane7_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane7_read_address1          ;
  wire                                          dma__memc__lane7_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane7_read_data1             ;
  wire                                          memc__dma__lane7_read_data_valid1       ;
  wire                                          memc__dma__lane7_read_ready1            ;
  wire                                          dma__memc__lane8_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane8_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane8_write_data1            ;
  wire                                          memc__dma__lane8_write_ready1           ;
  wire                                          dma__memc__lane8_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane8_read_address1          ;
  wire                                          dma__memc__lane8_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane8_read_data1             ;
  wire                                          memc__dma__lane8_read_data_valid1       ;
  wire                                          memc__dma__lane8_read_ready1            ;
  wire                                          dma__memc__lane9_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane9_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane9_write_data1            ;
  wire                                          memc__dma__lane9_write_ready1           ;
  wire                                          dma__memc__lane9_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane9_read_address1          ;
  wire                                          dma__memc__lane9_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane9_read_data1             ;
  wire                                          memc__dma__lane9_read_data_valid1       ;
  wire                                          memc__dma__lane9_read_ready1            ;
  wire                                          dma__memc__lane10_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane10_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane10_write_data1            ;
  wire                                          memc__dma__lane10_write_ready1           ;
  wire                                          dma__memc__lane10_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane10_read_address1          ;
  wire                                          dma__memc__lane10_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane10_read_data1             ;
  wire                                          memc__dma__lane10_read_data_valid1       ;
  wire                                          memc__dma__lane10_read_ready1            ;
  wire                                          dma__memc__lane11_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane11_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane11_write_data1            ;
  wire                                          memc__dma__lane11_write_ready1           ;
  wire                                          dma__memc__lane11_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane11_read_address1          ;
  wire                                          dma__memc__lane11_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane11_read_data1             ;
  wire                                          memc__dma__lane11_read_data_valid1       ;
  wire                                          memc__dma__lane11_read_ready1            ;
  wire                                          dma__memc__lane12_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane12_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane12_write_data1            ;
  wire                                          memc__dma__lane12_write_ready1           ;
  wire                                          dma__memc__lane12_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane12_read_address1          ;
  wire                                          dma__memc__lane12_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane12_read_data1             ;
  wire                                          memc__dma__lane12_read_data_valid1       ;
  wire                                          memc__dma__lane12_read_ready1            ;
  wire                                          dma__memc__lane13_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane13_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane13_write_data1            ;
  wire                                          memc__dma__lane13_write_ready1           ;
  wire                                          dma__memc__lane13_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane13_read_address1          ;
  wire                                          dma__memc__lane13_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane13_read_data1             ;
  wire                                          memc__dma__lane13_read_data_valid1       ;
  wire                                          memc__dma__lane13_read_ready1            ;
  wire                                          dma__memc__lane14_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane14_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane14_write_data1            ;
  wire                                          memc__dma__lane14_write_ready1           ;
  wire                                          dma__memc__lane14_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane14_read_address1          ;
  wire                                          dma__memc__lane14_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane14_read_data1             ;
  wire                                          memc__dma__lane14_read_data_valid1       ;
  wire                                          memc__dma__lane14_read_ready1            ;
  wire                                          dma__memc__lane15_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane15_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane15_write_data1            ;
  wire                                          memc__dma__lane15_write_ready1           ;
  wire                                          dma__memc__lane15_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane15_read_address1          ;
  wire                                          dma__memc__lane15_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane15_read_data1             ;
  wire                                          memc__dma__lane15_read_data_valid1       ;
  wire                                          memc__dma__lane15_read_ready1            ;
  wire                                          dma__memc__lane16_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane16_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane16_write_data1            ;
  wire                                          memc__dma__lane16_write_ready1           ;
  wire                                          dma__memc__lane16_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane16_read_address1          ;
  wire                                          dma__memc__lane16_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane16_read_data1             ;
  wire                                          memc__dma__lane16_read_data_valid1       ;
  wire                                          memc__dma__lane16_read_ready1            ;
  wire                                          dma__memc__lane17_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane17_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane17_write_data1            ;
  wire                                          memc__dma__lane17_write_ready1           ;
  wire                                          dma__memc__lane17_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane17_read_address1          ;
  wire                                          dma__memc__lane17_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane17_read_data1             ;
  wire                                          memc__dma__lane17_read_data_valid1       ;
  wire                                          memc__dma__lane17_read_ready1            ;
  wire                                          dma__memc__lane18_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane18_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane18_write_data1            ;
  wire                                          memc__dma__lane18_write_ready1           ;
  wire                                          dma__memc__lane18_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane18_read_address1          ;
  wire                                          dma__memc__lane18_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane18_read_data1             ;
  wire                                          memc__dma__lane18_read_data_valid1       ;
  wire                                          memc__dma__lane18_read_ready1            ;
  wire                                          dma__memc__lane19_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane19_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane19_write_data1            ;
  wire                                          memc__dma__lane19_write_ready1           ;
  wire                                          dma__memc__lane19_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane19_read_address1          ;
  wire                                          dma__memc__lane19_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane19_read_data1             ;
  wire                                          memc__dma__lane19_read_data_valid1       ;
  wire                                          memc__dma__lane19_read_ready1            ;
  wire                                          dma__memc__lane20_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane20_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane20_write_data1            ;
  wire                                          memc__dma__lane20_write_ready1           ;
  wire                                          dma__memc__lane20_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane20_read_address1          ;
  wire                                          dma__memc__lane20_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane20_read_data1             ;
  wire                                          memc__dma__lane20_read_data_valid1       ;
  wire                                          memc__dma__lane20_read_ready1            ;
  wire                                          dma__memc__lane21_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane21_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane21_write_data1            ;
  wire                                          memc__dma__lane21_write_ready1           ;
  wire                                          dma__memc__lane21_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane21_read_address1          ;
  wire                                          dma__memc__lane21_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane21_read_data1             ;
  wire                                          memc__dma__lane21_read_data_valid1       ;
  wire                                          memc__dma__lane21_read_ready1            ;
  wire                                          dma__memc__lane22_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane22_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane22_write_data1            ;
  wire                                          memc__dma__lane22_write_ready1           ;
  wire                                          dma__memc__lane22_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane22_read_address1          ;
  wire                                          dma__memc__lane22_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane22_read_data1             ;
  wire                                          memc__dma__lane22_read_data_valid1       ;
  wire                                          memc__dma__lane22_read_ready1            ;
  wire                                          dma__memc__lane23_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane23_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane23_write_data1            ;
  wire                                          memc__dma__lane23_write_ready1           ;
  wire                                          dma__memc__lane23_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane23_read_address1          ;
  wire                                          dma__memc__lane23_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane23_read_data1             ;
  wire                                          memc__dma__lane23_read_data_valid1       ;
  wire                                          memc__dma__lane23_read_ready1            ;
  wire                                          dma__memc__lane24_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane24_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane24_write_data1            ;
  wire                                          memc__dma__lane24_write_ready1           ;
  wire                                          dma__memc__lane24_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane24_read_address1          ;
  wire                                          dma__memc__lane24_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane24_read_data1             ;
  wire                                          memc__dma__lane24_read_data_valid1       ;
  wire                                          memc__dma__lane24_read_ready1            ;
  wire                                          dma__memc__lane25_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane25_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane25_write_data1            ;
  wire                                          memc__dma__lane25_write_ready1           ;
  wire                                          dma__memc__lane25_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane25_read_address1          ;
  wire                                          dma__memc__lane25_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane25_read_data1             ;
  wire                                          memc__dma__lane25_read_data_valid1       ;
  wire                                          memc__dma__lane25_read_ready1            ;
  wire                                          dma__memc__lane26_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane26_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane26_write_data1            ;
  wire                                          memc__dma__lane26_write_ready1           ;
  wire                                          dma__memc__lane26_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane26_read_address1          ;
  wire                                          dma__memc__lane26_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane26_read_data1             ;
  wire                                          memc__dma__lane26_read_data_valid1       ;
  wire                                          memc__dma__lane26_read_ready1            ;
  wire                                          dma__memc__lane27_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane27_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane27_write_data1            ;
  wire                                          memc__dma__lane27_write_ready1           ;
  wire                                          dma__memc__lane27_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane27_read_address1          ;
  wire                                          dma__memc__lane27_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane27_read_data1             ;
  wire                                          memc__dma__lane27_read_data_valid1       ;
  wire                                          memc__dma__lane27_read_ready1            ;
  wire                                          dma__memc__lane28_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane28_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane28_write_data1            ;
  wire                                          memc__dma__lane28_write_ready1           ;
  wire                                          dma__memc__lane28_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane28_read_address1          ;
  wire                                          dma__memc__lane28_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane28_read_data1             ;
  wire                                          memc__dma__lane28_read_data_valid1       ;
  wire                                          memc__dma__lane28_read_ready1            ;
  wire                                          dma__memc__lane29_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane29_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane29_write_data1            ;
  wire                                          memc__dma__lane29_write_ready1           ;
  wire                                          dma__memc__lane29_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane29_read_address1          ;
  wire                                          dma__memc__lane29_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane29_read_data1             ;
  wire                                          memc__dma__lane29_read_data_valid1       ;
  wire                                          memc__dma__lane29_read_ready1            ;
  wire                                          dma__memc__lane30_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane30_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane30_write_data1            ;
  wire                                          memc__dma__lane30_write_ready1           ;
  wire                                          dma__memc__lane30_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane30_read_address1          ;
  wire                                          dma__memc__lane30_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane30_read_data1             ;
  wire                                          memc__dma__lane30_read_data_valid1       ;
  wire                                          memc__dma__lane30_read_ready1            ;
  wire                                          dma__memc__lane31_write_valid1           ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane31_write_address1         ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  dma__memc__lane31_write_data1            ;
  wire                                          memc__dma__lane31_write_ready1           ;
  wire                                          dma__memc__lane31_read_valid1            ;
  wire   [`MEM_ACC_CONT_MEMORY_ADDRESS_RANGE ]  dma__memc__lane31_read_address1          ;
  wire                                          dma__memc__lane31_read_pause1            ;
  wire   [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__lane31_read_data1             ;
  wire                                          memc__dma__lane31_read_data_valid1       ;
  wire                                          memc__dma__lane31_read_ready1            ;

