
  // General control and status                                       
  assign    sys__pe0__allSynchronized     =    mgr0__sys__allSynchronized   ;
  assign    sys__mgr0__thisSynchronized   =    pe0__sys__thisSynchronized   ;
  assign    sys__mgr0__ready              =    pe0__sys__ready              ;
  assign    sys__mgr0__complete           =    pe0__sys__complete           ;

  // General control and status                                       
  assign    sys__pe1__allSynchronized     =    mgr1__sys__allSynchronized   ;
  assign    sys__mgr1__thisSynchronized   =    pe1__sys__thisSynchronized   ;
  assign    sys__mgr1__ready              =    pe1__sys__ready              ;
  assign    sys__mgr1__complete           =    pe1__sys__complete           ;

  // General control and status                                       
  assign    sys__pe2__allSynchronized     =    mgr2__sys__allSynchronized   ;
  assign    sys__mgr2__thisSynchronized   =    pe2__sys__thisSynchronized   ;
  assign    sys__mgr2__ready              =    pe2__sys__ready              ;
  assign    sys__mgr2__complete           =    pe2__sys__complete           ;

  // General control and status                                       
  assign    sys__pe3__allSynchronized     =    mgr3__sys__allSynchronized   ;
  assign    sys__mgr3__thisSynchronized   =    pe3__sys__thisSynchronized   ;
  assign    sys__mgr3__ready              =    pe3__sys__ready              ;
  assign    sys__mgr3__complete           =    pe3__sys__complete           ;

  // General control and status                                       
  assign    sys__pe4__allSynchronized     =    mgr4__sys__allSynchronized   ;
  assign    sys__mgr4__thisSynchronized   =    pe4__sys__thisSynchronized   ;
  assign    sys__mgr4__ready              =    pe4__sys__ready              ;
  assign    sys__mgr4__complete           =    pe4__sys__complete           ;

  // General control and status                                       
  assign    sys__pe5__allSynchronized     =    mgr5__sys__allSynchronized   ;
  assign    sys__mgr5__thisSynchronized   =    pe5__sys__thisSynchronized   ;
  assign    sys__mgr5__ready              =    pe5__sys__ready              ;
  assign    sys__mgr5__complete           =    pe5__sys__complete           ;

  // General control and status                                       
  assign    sys__pe6__allSynchronized     =    mgr6__sys__allSynchronized   ;
  assign    sys__mgr6__thisSynchronized   =    pe6__sys__thisSynchronized   ;
  assign    sys__mgr6__ready              =    pe6__sys__ready              ;
  assign    sys__mgr6__complete           =    pe6__sys__complete           ;

  // General control and status                                       
  assign    sys__pe7__allSynchronized     =    mgr7__sys__allSynchronized   ;
  assign    sys__mgr7__thisSynchronized   =    pe7__sys__thisSynchronized   ;
  assign    sys__mgr7__ready              =    pe7__sys__ready              ;
  assign    sys__mgr7__complete           =    pe7__sys__complete           ;

  // General control and status                                       
  assign    sys__pe8__allSynchronized     =    mgr8__sys__allSynchronized   ;
  assign    sys__mgr8__thisSynchronized   =    pe8__sys__thisSynchronized   ;
  assign    sys__mgr8__ready              =    pe8__sys__ready              ;
  assign    sys__mgr8__complete           =    pe8__sys__complete           ;

  // General control and status                                       
  assign    sys__pe9__allSynchronized     =    mgr9__sys__allSynchronized   ;
  assign    sys__mgr9__thisSynchronized   =    pe9__sys__thisSynchronized   ;
  assign    sys__mgr9__ready              =    pe9__sys__ready              ;
  assign    sys__mgr9__complete           =    pe9__sys__complete           ;

  // General control and status                                       
  assign    sys__pe10__allSynchronized     =    mgr10__sys__allSynchronized   ;
  assign    sys__mgr10__thisSynchronized   =    pe10__sys__thisSynchronized   ;
  assign    sys__mgr10__ready              =    pe10__sys__ready              ;
  assign    sys__mgr10__complete           =    pe10__sys__complete           ;

  // General control and status                                       
  assign    sys__pe11__allSynchronized     =    mgr11__sys__allSynchronized   ;
  assign    sys__mgr11__thisSynchronized   =    pe11__sys__thisSynchronized   ;
  assign    sys__mgr11__ready              =    pe11__sys__ready              ;
  assign    sys__mgr11__complete           =    pe11__sys__complete           ;

  // General control and status                                       
  assign    sys__pe12__allSynchronized     =    mgr12__sys__allSynchronized   ;
  assign    sys__mgr12__thisSynchronized   =    pe12__sys__thisSynchronized   ;
  assign    sys__mgr12__ready              =    pe12__sys__ready              ;
  assign    sys__mgr12__complete           =    pe12__sys__complete           ;

  // General control and status                                       
  assign    sys__pe13__allSynchronized     =    mgr13__sys__allSynchronized   ;
  assign    sys__mgr13__thisSynchronized   =    pe13__sys__thisSynchronized   ;
  assign    sys__mgr13__ready              =    pe13__sys__ready              ;
  assign    sys__mgr13__complete           =    pe13__sys__complete           ;

  // General control and status                                       
  assign    sys__pe14__allSynchronized     =    mgr14__sys__allSynchronized   ;
  assign    sys__mgr14__thisSynchronized   =    pe14__sys__thisSynchronized   ;
  assign    sys__mgr14__ready              =    pe14__sys__ready              ;
  assign    sys__mgr14__complete           =    pe14__sys__complete           ;

  // General control and status                                       
  assign    sys__pe15__allSynchronized     =    mgr15__sys__allSynchronized   ;
  assign    sys__mgr15__thisSynchronized   =    pe15__sys__thisSynchronized   ;
  assign    sys__mgr15__ready              =    pe15__sys__ready              ;
  assign    sys__mgr15__complete           =    pe15__sys__complete           ;

  // General control and status                                       
  assign    sys__pe16__allSynchronized     =    mgr16__sys__allSynchronized   ;
  assign    sys__mgr16__thisSynchronized   =    pe16__sys__thisSynchronized   ;
  assign    sys__mgr16__ready              =    pe16__sys__ready              ;
  assign    sys__mgr16__complete           =    pe16__sys__complete           ;

  // General control and status                                       
  assign    sys__pe17__allSynchronized     =    mgr17__sys__allSynchronized   ;
  assign    sys__mgr17__thisSynchronized   =    pe17__sys__thisSynchronized   ;
  assign    sys__mgr17__ready              =    pe17__sys__ready              ;
  assign    sys__mgr17__complete           =    pe17__sys__complete           ;

  // General control and status                                       
  assign    sys__pe18__allSynchronized     =    mgr18__sys__allSynchronized   ;
  assign    sys__mgr18__thisSynchronized   =    pe18__sys__thisSynchronized   ;
  assign    sys__mgr18__ready              =    pe18__sys__ready              ;
  assign    sys__mgr18__complete           =    pe18__sys__complete           ;

  // General control and status                                       
  assign    sys__pe19__allSynchronized     =    mgr19__sys__allSynchronized   ;
  assign    sys__mgr19__thisSynchronized   =    pe19__sys__thisSynchronized   ;
  assign    sys__mgr19__ready              =    pe19__sys__ready              ;
  assign    sys__mgr19__complete           =    pe19__sys__complete           ;

  // General control and status                                       
  assign    sys__pe20__allSynchronized     =    mgr20__sys__allSynchronized   ;
  assign    sys__mgr20__thisSynchronized   =    pe20__sys__thisSynchronized   ;
  assign    sys__mgr20__ready              =    pe20__sys__ready              ;
  assign    sys__mgr20__complete           =    pe20__sys__complete           ;

  // General control and status                                       
  assign    sys__pe21__allSynchronized     =    mgr21__sys__allSynchronized   ;
  assign    sys__mgr21__thisSynchronized   =    pe21__sys__thisSynchronized   ;
  assign    sys__mgr21__ready              =    pe21__sys__ready              ;
  assign    sys__mgr21__complete           =    pe21__sys__complete           ;

  // General control and status                                       
  assign    sys__pe22__allSynchronized     =    mgr22__sys__allSynchronized   ;
  assign    sys__mgr22__thisSynchronized   =    pe22__sys__thisSynchronized   ;
  assign    sys__mgr22__ready              =    pe22__sys__ready              ;
  assign    sys__mgr22__complete           =    pe22__sys__complete           ;

  // General control and status                                       
  assign    sys__pe23__allSynchronized     =    mgr23__sys__allSynchronized   ;
  assign    sys__mgr23__thisSynchronized   =    pe23__sys__thisSynchronized   ;
  assign    sys__mgr23__ready              =    pe23__sys__ready              ;
  assign    sys__mgr23__complete           =    pe23__sys__complete           ;

  // General control and status                                       
  assign    sys__pe24__allSynchronized     =    mgr24__sys__allSynchronized   ;
  assign    sys__mgr24__thisSynchronized   =    pe24__sys__thisSynchronized   ;
  assign    sys__mgr24__ready              =    pe24__sys__ready              ;
  assign    sys__mgr24__complete           =    pe24__sys__complete           ;

  // General control and status                                       
  assign    sys__pe25__allSynchronized     =    mgr25__sys__allSynchronized   ;
  assign    sys__mgr25__thisSynchronized   =    pe25__sys__thisSynchronized   ;
  assign    sys__mgr25__ready              =    pe25__sys__ready              ;
  assign    sys__mgr25__complete           =    pe25__sys__complete           ;

  // General control and status                                       
  assign    sys__pe26__allSynchronized     =    mgr26__sys__allSynchronized   ;
  assign    sys__mgr26__thisSynchronized   =    pe26__sys__thisSynchronized   ;
  assign    sys__mgr26__ready              =    pe26__sys__ready              ;
  assign    sys__mgr26__complete           =    pe26__sys__complete           ;

  // General control and status                                       
  assign    sys__pe27__allSynchronized     =    mgr27__sys__allSynchronized   ;
  assign    sys__mgr27__thisSynchronized   =    pe27__sys__thisSynchronized   ;
  assign    sys__mgr27__ready              =    pe27__sys__ready              ;
  assign    sys__mgr27__complete           =    pe27__sys__complete           ;

  // General control and status                                       
  assign    sys__pe28__allSynchronized     =    mgr28__sys__allSynchronized   ;
  assign    sys__mgr28__thisSynchronized   =    pe28__sys__thisSynchronized   ;
  assign    sys__mgr28__ready              =    pe28__sys__ready              ;
  assign    sys__mgr28__complete           =    pe28__sys__complete           ;

  // General control and status                                       
  assign    sys__pe29__allSynchronized     =    mgr29__sys__allSynchronized   ;
  assign    sys__mgr29__thisSynchronized   =    pe29__sys__thisSynchronized   ;
  assign    sys__mgr29__ready              =    pe29__sys__ready              ;
  assign    sys__mgr29__complete           =    pe29__sys__complete           ;

  // General control and status                                       
  assign    sys__pe30__allSynchronized     =    mgr30__sys__allSynchronized   ;
  assign    sys__mgr30__thisSynchronized   =    pe30__sys__thisSynchronized   ;
  assign    sys__mgr30__ready              =    pe30__sys__ready              ;
  assign    sys__mgr30__complete           =    pe30__sys__complete           ;

  // General control and status                                       
  assign    sys__pe31__allSynchronized     =    mgr31__sys__allSynchronized   ;
  assign    sys__mgr31__thisSynchronized   =    pe31__sys__thisSynchronized   ;
  assign    sys__mgr31__ready              =    pe31__sys__ready              ;
  assign    sys__mgr31__complete           =    pe31__sys__complete           ;

  // General control and status                                       
  assign    sys__pe32__allSynchronized     =    mgr32__sys__allSynchronized   ;
  assign    sys__mgr32__thisSynchronized   =    pe32__sys__thisSynchronized   ;
  assign    sys__mgr32__ready              =    pe32__sys__ready              ;
  assign    sys__mgr32__complete           =    pe32__sys__complete           ;

  // General control and status                                       
  assign    sys__pe33__allSynchronized     =    mgr33__sys__allSynchronized   ;
  assign    sys__mgr33__thisSynchronized   =    pe33__sys__thisSynchronized   ;
  assign    sys__mgr33__ready              =    pe33__sys__ready              ;
  assign    sys__mgr33__complete           =    pe33__sys__complete           ;

  // General control and status                                       
  assign    sys__pe34__allSynchronized     =    mgr34__sys__allSynchronized   ;
  assign    sys__mgr34__thisSynchronized   =    pe34__sys__thisSynchronized   ;
  assign    sys__mgr34__ready              =    pe34__sys__ready              ;
  assign    sys__mgr34__complete           =    pe34__sys__complete           ;

  // General control and status                                       
  assign    sys__pe35__allSynchronized     =    mgr35__sys__allSynchronized   ;
  assign    sys__mgr35__thisSynchronized   =    pe35__sys__thisSynchronized   ;
  assign    sys__mgr35__ready              =    pe35__sys__ready              ;
  assign    sys__mgr35__complete           =    pe35__sys__complete           ;

  // General control and status                                       
  assign    sys__pe36__allSynchronized     =    mgr36__sys__allSynchronized   ;
  assign    sys__mgr36__thisSynchronized   =    pe36__sys__thisSynchronized   ;
  assign    sys__mgr36__ready              =    pe36__sys__ready              ;
  assign    sys__mgr36__complete           =    pe36__sys__complete           ;

  // General control and status                                       
  assign    sys__pe37__allSynchronized     =    mgr37__sys__allSynchronized   ;
  assign    sys__mgr37__thisSynchronized   =    pe37__sys__thisSynchronized   ;
  assign    sys__mgr37__ready              =    pe37__sys__ready              ;
  assign    sys__mgr37__complete           =    pe37__sys__complete           ;

  // General control and status                                       
  assign    sys__pe38__allSynchronized     =    mgr38__sys__allSynchronized   ;
  assign    sys__mgr38__thisSynchronized   =    pe38__sys__thisSynchronized   ;
  assign    sys__mgr38__ready              =    pe38__sys__ready              ;
  assign    sys__mgr38__complete           =    pe38__sys__complete           ;

  // General control and status                                       
  assign    sys__pe39__allSynchronized     =    mgr39__sys__allSynchronized   ;
  assign    sys__mgr39__thisSynchronized   =    pe39__sys__thisSynchronized   ;
  assign    sys__mgr39__ready              =    pe39__sys__ready              ;
  assign    sys__mgr39__complete           =    pe39__sys__complete           ;

  // General control and status                                       
  assign    sys__pe40__allSynchronized     =    mgr40__sys__allSynchronized   ;
  assign    sys__mgr40__thisSynchronized   =    pe40__sys__thisSynchronized   ;
  assign    sys__mgr40__ready              =    pe40__sys__ready              ;
  assign    sys__mgr40__complete           =    pe40__sys__complete           ;

  // General control and status                                       
  assign    sys__pe41__allSynchronized     =    mgr41__sys__allSynchronized   ;
  assign    sys__mgr41__thisSynchronized   =    pe41__sys__thisSynchronized   ;
  assign    sys__mgr41__ready              =    pe41__sys__ready              ;
  assign    sys__mgr41__complete           =    pe41__sys__complete           ;

  // General control and status                                       
  assign    sys__pe42__allSynchronized     =    mgr42__sys__allSynchronized   ;
  assign    sys__mgr42__thisSynchronized   =    pe42__sys__thisSynchronized   ;
  assign    sys__mgr42__ready              =    pe42__sys__ready              ;
  assign    sys__mgr42__complete           =    pe42__sys__complete           ;

  // General control and status                                       
  assign    sys__pe43__allSynchronized     =    mgr43__sys__allSynchronized   ;
  assign    sys__mgr43__thisSynchronized   =    pe43__sys__thisSynchronized   ;
  assign    sys__mgr43__ready              =    pe43__sys__ready              ;
  assign    sys__mgr43__complete           =    pe43__sys__complete           ;

  // General control and status                                       
  assign    sys__pe44__allSynchronized     =    mgr44__sys__allSynchronized   ;
  assign    sys__mgr44__thisSynchronized   =    pe44__sys__thisSynchronized   ;
  assign    sys__mgr44__ready              =    pe44__sys__ready              ;
  assign    sys__mgr44__complete           =    pe44__sys__complete           ;

  // General control and status                                       
  assign    sys__pe45__allSynchronized     =    mgr45__sys__allSynchronized   ;
  assign    sys__mgr45__thisSynchronized   =    pe45__sys__thisSynchronized   ;
  assign    sys__mgr45__ready              =    pe45__sys__ready              ;
  assign    sys__mgr45__complete           =    pe45__sys__complete           ;

  // General control and status                                       
  assign    sys__pe46__allSynchronized     =    mgr46__sys__allSynchronized   ;
  assign    sys__mgr46__thisSynchronized   =    pe46__sys__thisSynchronized   ;
  assign    sys__mgr46__ready              =    pe46__sys__ready              ;
  assign    sys__mgr46__complete           =    pe46__sys__complete           ;

  // General control and status                                       
  assign    sys__pe47__allSynchronized     =    mgr47__sys__allSynchronized   ;
  assign    sys__mgr47__thisSynchronized   =    pe47__sys__thisSynchronized   ;
  assign    sys__mgr47__ready              =    pe47__sys__ready              ;
  assign    sys__mgr47__complete           =    pe47__sys__complete           ;

  // General control and status                                       
  assign    sys__pe48__allSynchronized     =    mgr48__sys__allSynchronized   ;
  assign    sys__mgr48__thisSynchronized   =    pe48__sys__thisSynchronized   ;
  assign    sys__mgr48__ready              =    pe48__sys__ready              ;
  assign    sys__mgr48__complete           =    pe48__sys__complete           ;

  // General control and status                                       
  assign    sys__pe49__allSynchronized     =    mgr49__sys__allSynchronized   ;
  assign    sys__mgr49__thisSynchronized   =    pe49__sys__thisSynchronized   ;
  assign    sys__mgr49__ready              =    pe49__sys__ready              ;
  assign    sys__mgr49__complete           =    pe49__sys__complete           ;

  // General control and status                                       
  assign    sys__pe50__allSynchronized     =    mgr50__sys__allSynchronized   ;
  assign    sys__mgr50__thisSynchronized   =    pe50__sys__thisSynchronized   ;
  assign    sys__mgr50__ready              =    pe50__sys__ready              ;
  assign    sys__mgr50__complete           =    pe50__sys__complete           ;

  // General control and status                                       
  assign    sys__pe51__allSynchronized     =    mgr51__sys__allSynchronized   ;
  assign    sys__mgr51__thisSynchronized   =    pe51__sys__thisSynchronized   ;
  assign    sys__mgr51__ready              =    pe51__sys__ready              ;
  assign    sys__mgr51__complete           =    pe51__sys__complete           ;

  // General control and status                                       
  assign    sys__pe52__allSynchronized     =    mgr52__sys__allSynchronized   ;
  assign    sys__mgr52__thisSynchronized   =    pe52__sys__thisSynchronized   ;
  assign    sys__mgr52__ready              =    pe52__sys__ready              ;
  assign    sys__mgr52__complete           =    pe52__sys__complete           ;

  // General control and status                                       
  assign    sys__pe53__allSynchronized     =    mgr53__sys__allSynchronized   ;
  assign    sys__mgr53__thisSynchronized   =    pe53__sys__thisSynchronized   ;
  assign    sys__mgr53__ready              =    pe53__sys__ready              ;
  assign    sys__mgr53__complete           =    pe53__sys__complete           ;

  // General control and status                                       
  assign    sys__pe54__allSynchronized     =    mgr54__sys__allSynchronized   ;
  assign    sys__mgr54__thisSynchronized   =    pe54__sys__thisSynchronized   ;
  assign    sys__mgr54__ready              =    pe54__sys__ready              ;
  assign    sys__mgr54__complete           =    pe54__sys__complete           ;

  // General control and status                                       
  assign    sys__pe55__allSynchronized     =    mgr55__sys__allSynchronized   ;
  assign    sys__mgr55__thisSynchronized   =    pe55__sys__thisSynchronized   ;
  assign    sys__mgr55__ready              =    pe55__sys__ready              ;
  assign    sys__mgr55__complete           =    pe55__sys__complete           ;

  // General control and status                                       
  assign    sys__pe56__allSynchronized     =    mgr56__sys__allSynchronized   ;
  assign    sys__mgr56__thisSynchronized   =    pe56__sys__thisSynchronized   ;
  assign    sys__mgr56__ready              =    pe56__sys__ready              ;
  assign    sys__mgr56__complete           =    pe56__sys__complete           ;

  // General control and status                                       
  assign    sys__pe57__allSynchronized     =    mgr57__sys__allSynchronized   ;
  assign    sys__mgr57__thisSynchronized   =    pe57__sys__thisSynchronized   ;
  assign    sys__mgr57__ready              =    pe57__sys__ready              ;
  assign    sys__mgr57__complete           =    pe57__sys__complete           ;

  // General control and status                                       
  assign    sys__pe58__allSynchronized     =    mgr58__sys__allSynchronized   ;
  assign    sys__mgr58__thisSynchronized   =    pe58__sys__thisSynchronized   ;
  assign    sys__mgr58__ready              =    pe58__sys__ready              ;
  assign    sys__mgr58__complete           =    pe58__sys__complete           ;

  // General control and status                                       
  assign    sys__pe59__allSynchronized     =    mgr59__sys__allSynchronized   ;
  assign    sys__mgr59__thisSynchronized   =    pe59__sys__thisSynchronized   ;
  assign    sys__mgr59__ready              =    pe59__sys__ready              ;
  assign    sys__mgr59__complete           =    pe59__sys__complete           ;

  // General control and status                                       
  assign    sys__pe60__allSynchronized     =    mgr60__sys__allSynchronized   ;
  assign    sys__mgr60__thisSynchronized   =    pe60__sys__thisSynchronized   ;
  assign    sys__mgr60__ready              =    pe60__sys__ready              ;
  assign    sys__mgr60__complete           =    pe60__sys__complete           ;

  // General control and status                                       
  assign    sys__pe61__allSynchronized     =    mgr61__sys__allSynchronized   ;
  assign    sys__mgr61__thisSynchronized   =    pe61__sys__thisSynchronized   ;
  assign    sys__mgr61__ready              =    pe61__sys__ready              ;
  assign    sys__mgr61__complete           =    pe61__sys__complete           ;

  // General control and status                                       
  assign    sys__pe62__allSynchronized     =    mgr62__sys__allSynchronized   ;
  assign    sys__mgr62__thisSynchronized   =    pe62__sys__thisSynchronized   ;
  assign    sys__mgr62__ready              =    pe62__sys__ready              ;
  assign    sys__mgr62__complete           =    pe62__sys__complete           ;

  // General control and status                                       
  assign    sys__pe63__allSynchronized     =    mgr63__sys__allSynchronized   ;
  assign    sys__mgr63__thisSynchronized   =    pe63__sys__thisSynchronized   ;
  assign    sys__mgr63__ready              =    pe63__sys__ready              ;
  assign    sys__mgr63__complete           =    pe63__sys__complete           ;
