
               // OOB carries PE configuration                                               
               .std__pe__oob_cntl                  ( std__pe__oob_cntl               ),      
               .std__pe__oob_valid                 ( std__pe__oob_valid              ),      
               .pe__std__oob_ready                 ( pe__std__oob_ready              ),      
               .std__pe__oob_type                  ( std__pe__oob_type               ),      
               .std__pe__oob_data                  ( std__pe__oob_data               ),      
