
  // Send an 'all' synchronized to all Managers's 
  // sys__mgr__thisSyncnronized basically means all the streams in a PE are complete
  // The PE controller will move to a 'final' state once it receives sys__pe__allSynchronized
  wire  mgr__sys__allSynchronized = mgr_inst[0].sys__mgr__thisSynchronized & 
                                   mgr_inst[1].sys__mgr__thisSynchronized & 
                                   mgr_inst[2].sys__mgr__thisSynchronized & 
                                   mgr_inst[3].sys__mgr__thisSynchronized & 
                                   mgr_inst[4].sys__mgr__thisSynchronized & 
                                   mgr_inst[5].sys__mgr__thisSynchronized & 
                                   mgr_inst[6].sys__mgr__thisSynchronized & 
                                   mgr_inst[7].sys__mgr__thisSynchronized & 
                                   mgr_inst[8].sys__mgr__thisSynchronized & 
                                   mgr_inst[9].sys__mgr__thisSynchronized & 
                                   mgr_inst[10].sys__mgr__thisSynchronized & 
                                   mgr_inst[11].sys__mgr__thisSynchronized & 
                                   mgr_inst[12].sys__mgr__thisSynchronized & 
                                   mgr_inst[13].sys__mgr__thisSynchronized & 
                                   mgr_inst[14].sys__mgr__thisSynchronized & 
                                   mgr_inst[15].sys__mgr__thisSynchronized & 
                                   mgr_inst[16].sys__mgr__thisSynchronized & 
                                   mgr_inst[17].sys__mgr__thisSynchronized & 
                                   mgr_inst[18].sys__mgr__thisSynchronized & 
                                   mgr_inst[19].sys__mgr__thisSynchronized & 
                                   mgr_inst[20].sys__mgr__thisSynchronized & 
                                   mgr_inst[21].sys__mgr__thisSynchronized & 
                                   mgr_inst[22].sys__mgr__thisSynchronized & 
                                   mgr_inst[23].sys__mgr__thisSynchronized & 
                                   mgr_inst[24].sys__mgr__thisSynchronized & 
                                   mgr_inst[25].sys__mgr__thisSynchronized & 
                                   mgr_inst[26].sys__mgr__thisSynchronized & 
                                   mgr_inst[27].sys__mgr__thisSynchronized & 
                                   mgr_inst[28].sys__mgr__thisSynchronized & 
                                   mgr_inst[29].sys__mgr__thisSynchronized & 
                                   mgr_inst[30].sys__mgr__thisSynchronized & 
                                   mgr_inst[31].sys__mgr__thisSynchronized & 
                                   mgr_inst[32].sys__mgr__thisSynchronized & 
                                   mgr_inst[33].sys__mgr__thisSynchronized & 
                                   mgr_inst[34].sys__mgr__thisSynchronized & 
                                   mgr_inst[35].sys__mgr__thisSynchronized & 
                                   mgr_inst[36].sys__mgr__thisSynchronized & 
                                   mgr_inst[37].sys__mgr__thisSynchronized & 
                                   mgr_inst[38].sys__mgr__thisSynchronized & 
                                   mgr_inst[39].sys__mgr__thisSynchronized & 
                                   mgr_inst[40].sys__mgr__thisSynchronized & 
                                   mgr_inst[41].sys__mgr__thisSynchronized & 
                                   mgr_inst[42].sys__mgr__thisSynchronized & 
                                   mgr_inst[43].sys__mgr__thisSynchronized & 
                                   mgr_inst[44].sys__mgr__thisSynchronized & 
                                   mgr_inst[45].sys__mgr__thisSynchronized & 
                                   mgr_inst[46].sys__mgr__thisSynchronized & 
                                   mgr_inst[47].sys__mgr__thisSynchronized & 
                                   mgr_inst[48].sys__mgr__thisSynchronized & 
                                   mgr_inst[49].sys__mgr__thisSynchronized & 
                                   mgr_inst[50].sys__mgr__thisSynchronized & 
                                   mgr_inst[51].sys__mgr__thisSynchronized & 
                                   mgr_inst[52].sys__mgr__thisSynchronized & 
                                   mgr_inst[53].sys__mgr__thisSynchronized & 
                                   mgr_inst[54].sys__mgr__thisSynchronized & 
                                   mgr_inst[55].sys__mgr__thisSynchronized & 
                                   mgr_inst[56].sys__mgr__thisSynchronized & 
                                   mgr_inst[57].sys__mgr__thisSynchronized & 
                                   mgr_inst[58].sys__mgr__thisSynchronized & 
                                   mgr_inst[59].sys__mgr__thisSynchronized & 
                                   mgr_inst[60].sys__mgr__thisSynchronized & 
                                   mgr_inst[61].sys__mgr__thisSynchronized & 
                                   mgr_inst[62].sys__mgr__thisSynchronized & 
                                   mgr_inst[63].sys__mgr__thisSynchronized ; 