
               // Lane 0                 
               .std__mgr__lane0_strm0_ready         ( std__mgr__lane0_strm0_ready      ),      
               .mgr__std__lane0_strm0_cntl          ( mgr__std__lane0_strm0_cntl       ),      
               .mgr__std__lane0_strm0_data          ( mgr__std__lane0_strm0_data       ),      
               .mgr__std__lane0_strm0_data_valid    ( mgr__std__lane0_strm0_data_valid ),      
               .std__mgr__lane0_strm1_ready         ( std__mgr__lane0_strm1_ready      ),      
               .mgr__std__lane0_strm1_cntl          ( mgr__std__lane0_strm1_cntl       ),      
               .mgr__std__lane0_strm1_data          ( mgr__std__lane0_strm1_data       ),      
               .mgr__std__lane0_strm1_data_valid    ( mgr__std__lane0_strm1_data_valid ),      
               // Lane 1                 
               .std__mgr__lane1_strm0_ready         ( std__mgr__lane1_strm0_ready      ),      
               .mgr__std__lane1_strm0_cntl          ( mgr__std__lane1_strm0_cntl       ),      
               .mgr__std__lane1_strm0_data          ( mgr__std__lane1_strm0_data       ),      
               .mgr__std__lane1_strm0_data_valid    ( mgr__std__lane1_strm0_data_valid ),      
               .std__mgr__lane1_strm1_ready         ( std__mgr__lane1_strm1_ready      ),      
               .mgr__std__lane1_strm1_cntl          ( mgr__std__lane1_strm1_cntl       ),      
               .mgr__std__lane1_strm1_data          ( mgr__std__lane1_strm1_data       ),      
               .mgr__std__lane1_strm1_data_valid    ( mgr__std__lane1_strm1_data_valid ),      
               // Lane 2                 
               .std__mgr__lane2_strm0_ready         ( std__mgr__lane2_strm0_ready      ),      
               .mgr__std__lane2_strm0_cntl          ( mgr__std__lane2_strm0_cntl       ),      
               .mgr__std__lane2_strm0_data          ( mgr__std__lane2_strm0_data       ),      
               .mgr__std__lane2_strm0_data_valid    ( mgr__std__lane2_strm0_data_valid ),      
               .std__mgr__lane2_strm1_ready         ( std__mgr__lane2_strm1_ready      ),      
               .mgr__std__lane2_strm1_cntl          ( mgr__std__lane2_strm1_cntl       ),      
               .mgr__std__lane2_strm1_data          ( mgr__std__lane2_strm1_data       ),      
               .mgr__std__lane2_strm1_data_valid    ( mgr__std__lane2_strm1_data_valid ),      
               // Lane 3                 
               .std__mgr__lane3_strm0_ready         ( std__mgr__lane3_strm0_ready      ),      
               .mgr__std__lane3_strm0_cntl          ( mgr__std__lane3_strm0_cntl       ),      
               .mgr__std__lane3_strm0_data          ( mgr__std__lane3_strm0_data       ),      
               .mgr__std__lane3_strm0_data_valid    ( mgr__std__lane3_strm0_data_valid ),      
               .std__mgr__lane3_strm1_ready         ( std__mgr__lane3_strm1_ready      ),      
               .mgr__std__lane3_strm1_cntl          ( mgr__std__lane3_strm1_cntl       ),      
               .mgr__std__lane3_strm1_data          ( mgr__std__lane3_strm1_data       ),      
               .mgr__std__lane3_strm1_data_valid    ( mgr__std__lane3_strm1_data_valid ),      
               // Lane 4                 
               .std__mgr__lane4_strm0_ready         ( std__mgr__lane4_strm0_ready      ),      
               .mgr__std__lane4_strm0_cntl          ( mgr__std__lane4_strm0_cntl       ),      
               .mgr__std__lane4_strm0_data          ( mgr__std__lane4_strm0_data       ),      
               .mgr__std__lane4_strm0_data_valid    ( mgr__std__lane4_strm0_data_valid ),      
               .std__mgr__lane4_strm1_ready         ( std__mgr__lane4_strm1_ready      ),      
               .mgr__std__lane4_strm1_cntl          ( mgr__std__lane4_strm1_cntl       ),      
               .mgr__std__lane4_strm1_data          ( mgr__std__lane4_strm1_data       ),      
               .mgr__std__lane4_strm1_data_valid    ( mgr__std__lane4_strm1_data_valid ),      
               // Lane 5                 
               .std__mgr__lane5_strm0_ready         ( std__mgr__lane5_strm0_ready      ),      
               .mgr__std__lane5_strm0_cntl          ( mgr__std__lane5_strm0_cntl       ),      
               .mgr__std__lane5_strm0_data          ( mgr__std__lane5_strm0_data       ),      
               .mgr__std__lane5_strm0_data_valid    ( mgr__std__lane5_strm0_data_valid ),      
               .std__mgr__lane5_strm1_ready         ( std__mgr__lane5_strm1_ready      ),      
               .mgr__std__lane5_strm1_cntl          ( mgr__std__lane5_strm1_cntl       ),      
               .mgr__std__lane5_strm1_data          ( mgr__std__lane5_strm1_data       ),      
               .mgr__std__lane5_strm1_data_valid    ( mgr__std__lane5_strm1_data_valid ),      
               // Lane 6                 
               .std__mgr__lane6_strm0_ready         ( std__mgr__lane6_strm0_ready      ),      
               .mgr__std__lane6_strm0_cntl          ( mgr__std__lane6_strm0_cntl       ),      
               .mgr__std__lane6_strm0_data          ( mgr__std__lane6_strm0_data       ),      
               .mgr__std__lane6_strm0_data_valid    ( mgr__std__lane6_strm0_data_valid ),      
               .std__mgr__lane6_strm1_ready         ( std__mgr__lane6_strm1_ready      ),      
               .mgr__std__lane6_strm1_cntl          ( mgr__std__lane6_strm1_cntl       ),      
               .mgr__std__lane6_strm1_data          ( mgr__std__lane6_strm1_data       ),      
               .mgr__std__lane6_strm1_data_valid    ( mgr__std__lane6_strm1_data_valid ),      
               // Lane 7                 
               .std__mgr__lane7_strm0_ready         ( std__mgr__lane7_strm0_ready      ),      
               .mgr__std__lane7_strm0_cntl          ( mgr__std__lane7_strm0_cntl       ),      
               .mgr__std__lane7_strm0_data          ( mgr__std__lane7_strm0_data       ),      
               .mgr__std__lane7_strm0_data_valid    ( mgr__std__lane7_strm0_data_valid ),      
               .std__mgr__lane7_strm1_ready         ( std__mgr__lane7_strm1_ready      ),      
               .mgr__std__lane7_strm1_cntl          ( mgr__std__lane7_strm1_cntl       ),      
               .mgr__std__lane7_strm1_data          ( mgr__std__lane7_strm1_data       ),      
               .mgr__std__lane7_strm1_data_valid    ( mgr__std__lane7_strm1_data_valid ),      
               // Lane 8                 
               .std__mgr__lane8_strm0_ready         ( std__mgr__lane8_strm0_ready      ),      
               .mgr__std__lane8_strm0_cntl          ( mgr__std__lane8_strm0_cntl       ),      
               .mgr__std__lane8_strm0_data          ( mgr__std__lane8_strm0_data       ),      
               .mgr__std__lane8_strm0_data_valid    ( mgr__std__lane8_strm0_data_valid ),      
               .std__mgr__lane8_strm1_ready         ( std__mgr__lane8_strm1_ready      ),      
               .mgr__std__lane8_strm1_cntl          ( mgr__std__lane8_strm1_cntl       ),      
               .mgr__std__lane8_strm1_data          ( mgr__std__lane8_strm1_data       ),      
               .mgr__std__lane8_strm1_data_valid    ( mgr__std__lane8_strm1_data_valid ),      
               // Lane 9                 
               .std__mgr__lane9_strm0_ready         ( std__mgr__lane9_strm0_ready      ),      
               .mgr__std__lane9_strm0_cntl          ( mgr__std__lane9_strm0_cntl       ),      
               .mgr__std__lane9_strm0_data          ( mgr__std__lane9_strm0_data       ),      
               .mgr__std__lane9_strm0_data_valid    ( mgr__std__lane9_strm0_data_valid ),      
               .std__mgr__lane9_strm1_ready         ( std__mgr__lane9_strm1_ready      ),      
               .mgr__std__lane9_strm1_cntl          ( mgr__std__lane9_strm1_cntl       ),      
               .mgr__std__lane9_strm1_data          ( mgr__std__lane9_strm1_data       ),      
               .mgr__std__lane9_strm1_data_valid    ( mgr__std__lane9_strm1_data_valid ),      
               // Lane 10                 
               .std__mgr__lane10_strm0_ready         ( std__mgr__lane10_strm0_ready      ),      
               .mgr__std__lane10_strm0_cntl          ( mgr__std__lane10_strm0_cntl       ),      
               .mgr__std__lane10_strm0_data          ( mgr__std__lane10_strm0_data       ),      
               .mgr__std__lane10_strm0_data_valid    ( mgr__std__lane10_strm0_data_valid ),      
               .std__mgr__lane10_strm1_ready         ( std__mgr__lane10_strm1_ready      ),      
               .mgr__std__lane10_strm1_cntl          ( mgr__std__lane10_strm1_cntl       ),      
               .mgr__std__lane10_strm1_data          ( mgr__std__lane10_strm1_data       ),      
               .mgr__std__lane10_strm1_data_valid    ( mgr__std__lane10_strm1_data_valid ),      
               // Lane 11                 
               .std__mgr__lane11_strm0_ready         ( std__mgr__lane11_strm0_ready      ),      
               .mgr__std__lane11_strm0_cntl          ( mgr__std__lane11_strm0_cntl       ),      
               .mgr__std__lane11_strm0_data          ( mgr__std__lane11_strm0_data       ),      
               .mgr__std__lane11_strm0_data_valid    ( mgr__std__lane11_strm0_data_valid ),      
               .std__mgr__lane11_strm1_ready         ( std__mgr__lane11_strm1_ready      ),      
               .mgr__std__lane11_strm1_cntl          ( mgr__std__lane11_strm1_cntl       ),      
               .mgr__std__lane11_strm1_data          ( mgr__std__lane11_strm1_data       ),      
               .mgr__std__lane11_strm1_data_valid    ( mgr__std__lane11_strm1_data_valid ),      
               // Lane 12                 
               .std__mgr__lane12_strm0_ready         ( std__mgr__lane12_strm0_ready      ),      
               .mgr__std__lane12_strm0_cntl          ( mgr__std__lane12_strm0_cntl       ),      
               .mgr__std__lane12_strm0_data          ( mgr__std__lane12_strm0_data       ),      
               .mgr__std__lane12_strm0_data_valid    ( mgr__std__lane12_strm0_data_valid ),      
               .std__mgr__lane12_strm1_ready         ( std__mgr__lane12_strm1_ready      ),      
               .mgr__std__lane12_strm1_cntl          ( mgr__std__lane12_strm1_cntl       ),      
               .mgr__std__lane12_strm1_data          ( mgr__std__lane12_strm1_data       ),      
               .mgr__std__lane12_strm1_data_valid    ( mgr__std__lane12_strm1_data_valid ),      
               // Lane 13                 
               .std__mgr__lane13_strm0_ready         ( std__mgr__lane13_strm0_ready      ),      
               .mgr__std__lane13_strm0_cntl          ( mgr__std__lane13_strm0_cntl       ),      
               .mgr__std__lane13_strm0_data          ( mgr__std__lane13_strm0_data       ),      
               .mgr__std__lane13_strm0_data_valid    ( mgr__std__lane13_strm0_data_valid ),      
               .std__mgr__lane13_strm1_ready         ( std__mgr__lane13_strm1_ready      ),      
               .mgr__std__lane13_strm1_cntl          ( mgr__std__lane13_strm1_cntl       ),      
               .mgr__std__lane13_strm1_data          ( mgr__std__lane13_strm1_data       ),      
               .mgr__std__lane13_strm1_data_valid    ( mgr__std__lane13_strm1_data_valid ),      
               // Lane 14                 
               .std__mgr__lane14_strm0_ready         ( std__mgr__lane14_strm0_ready      ),      
               .mgr__std__lane14_strm0_cntl          ( mgr__std__lane14_strm0_cntl       ),      
               .mgr__std__lane14_strm0_data          ( mgr__std__lane14_strm0_data       ),      
               .mgr__std__lane14_strm0_data_valid    ( mgr__std__lane14_strm0_data_valid ),      
               .std__mgr__lane14_strm1_ready         ( std__mgr__lane14_strm1_ready      ),      
               .mgr__std__lane14_strm1_cntl          ( mgr__std__lane14_strm1_cntl       ),      
               .mgr__std__lane14_strm1_data          ( mgr__std__lane14_strm1_data       ),      
               .mgr__std__lane14_strm1_data_valid    ( mgr__std__lane14_strm1_data_valid ),      
               // Lane 15                 
               .std__mgr__lane15_strm0_ready         ( std__mgr__lane15_strm0_ready      ),      
               .mgr__std__lane15_strm0_cntl          ( mgr__std__lane15_strm0_cntl       ),      
               .mgr__std__lane15_strm0_data          ( mgr__std__lane15_strm0_data       ),      
               .mgr__std__lane15_strm0_data_valid    ( mgr__std__lane15_strm0_data_valid ),      
               .std__mgr__lane15_strm1_ready         ( std__mgr__lane15_strm1_ready      ),      
               .mgr__std__lane15_strm1_cntl          ( mgr__std__lane15_strm1_cntl       ),      
               .mgr__std__lane15_strm1_data          ( mgr__std__lane15_strm1_data       ),      
               .mgr__std__lane15_strm1_data_valid    ( mgr__std__lane15_strm1_data_valid ),      
               // Lane 16                 
               .std__mgr__lane16_strm0_ready         ( std__mgr__lane16_strm0_ready      ),      
               .mgr__std__lane16_strm0_cntl          ( mgr__std__lane16_strm0_cntl       ),      
               .mgr__std__lane16_strm0_data          ( mgr__std__lane16_strm0_data       ),      
               .mgr__std__lane16_strm0_data_valid    ( mgr__std__lane16_strm0_data_valid ),      
               .std__mgr__lane16_strm1_ready         ( std__mgr__lane16_strm1_ready      ),      
               .mgr__std__lane16_strm1_cntl          ( mgr__std__lane16_strm1_cntl       ),      
               .mgr__std__lane16_strm1_data          ( mgr__std__lane16_strm1_data       ),      
               .mgr__std__lane16_strm1_data_valid    ( mgr__std__lane16_strm1_data_valid ),      
               // Lane 17                 
               .std__mgr__lane17_strm0_ready         ( std__mgr__lane17_strm0_ready      ),      
               .mgr__std__lane17_strm0_cntl          ( mgr__std__lane17_strm0_cntl       ),      
               .mgr__std__lane17_strm0_data          ( mgr__std__lane17_strm0_data       ),      
               .mgr__std__lane17_strm0_data_valid    ( mgr__std__lane17_strm0_data_valid ),      
               .std__mgr__lane17_strm1_ready         ( std__mgr__lane17_strm1_ready      ),      
               .mgr__std__lane17_strm1_cntl          ( mgr__std__lane17_strm1_cntl       ),      
               .mgr__std__lane17_strm1_data          ( mgr__std__lane17_strm1_data       ),      
               .mgr__std__lane17_strm1_data_valid    ( mgr__std__lane17_strm1_data_valid ),      
               // Lane 18                 
               .std__mgr__lane18_strm0_ready         ( std__mgr__lane18_strm0_ready      ),      
               .mgr__std__lane18_strm0_cntl          ( mgr__std__lane18_strm0_cntl       ),      
               .mgr__std__lane18_strm0_data          ( mgr__std__lane18_strm0_data       ),      
               .mgr__std__lane18_strm0_data_valid    ( mgr__std__lane18_strm0_data_valid ),      
               .std__mgr__lane18_strm1_ready         ( std__mgr__lane18_strm1_ready      ),      
               .mgr__std__lane18_strm1_cntl          ( mgr__std__lane18_strm1_cntl       ),      
               .mgr__std__lane18_strm1_data          ( mgr__std__lane18_strm1_data       ),      
               .mgr__std__lane18_strm1_data_valid    ( mgr__std__lane18_strm1_data_valid ),      
               // Lane 19                 
               .std__mgr__lane19_strm0_ready         ( std__mgr__lane19_strm0_ready      ),      
               .mgr__std__lane19_strm0_cntl          ( mgr__std__lane19_strm0_cntl       ),      
               .mgr__std__lane19_strm0_data          ( mgr__std__lane19_strm0_data       ),      
               .mgr__std__lane19_strm0_data_valid    ( mgr__std__lane19_strm0_data_valid ),      
               .std__mgr__lane19_strm1_ready         ( std__mgr__lane19_strm1_ready      ),      
               .mgr__std__lane19_strm1_cntl          ( mgr__std__lane19_strm1_cntl       ),      
               .mgr__std__lane19_strm1_data          ( mgr__std__lane19_strm1_data       ),      
               .mgr__std__lane19_strm1_data_valid    ( mgr__std__lane19_strm1_data_valid ),      
               // Lane 20                 
               .std__mgr__lane20_strm0_ready         ( std__mgr__lane20_strm0_ready      ),      
               .mgr__std__lane20_strm0_cntl          ( mgr__std__lane20_strm0_cntl       ),      
               .mgr__std__lane20_strm0_data          ( mgr__std__lane20_strm0_data       ),      
               .mgr__std__lane20_strm0_data_valid    ( mgr__std__lane20_strm0_data_valid ),      
               .std__mgr__lane20_strm1_ready         ( std__mgr__lane20_strm1_ready      ),      
               .mgr__std__lane20_strm1_cntl          ( mgr__std__lane20_strm1_cntl       ),      
               .mgr__std__lane20_strm1_data          ( mgr__std__lane20_strm1_data       ),      
               .mgr__std__lane20_strm1_data_valid    ( mgr__std__lane20_strm1_data_valid ),      
               // Lane 21                 
               .std__mgr__lane21_strm0_ready         ( std__mgr__lane21_strm0_ready      ),      
               .mgr__std__lane21_strm0_cntl          ( mgr__std__lane21_strm0_cntl       ),      
               .mgr__std__lane21_strm0_data          ( mgr__std__lane21_strm0_data       ),      
               .mgr__std__lane21_strm0_data_valid    ( mgr__std__lane21_strm0_data_valid ),      
               .std__mgr__lane21_strm1_ready         ( std__mgr__lane21_strm1_ready      ),      
               .mgr__std__lane21_strm1_cntl          ( mgr__std__lane21_strm1_cntl       ),      
               .mgr__std__lane21_strm1_data          ( mgr__std__lane21_strm1_data       ),      
               .mgr__std__lane21_strm1_data_valid    ( mgr__std__lane21_strm1_data_valid ),      
               // Lane 22                 
               .std__mgr__lane22_strm0_ready         ( std__mgr__lane22_strm0_ready      ),      
               .mgr__std__lane22_strm0_cntl          ( mgr__std__lane22_strm0_cntl       ),      
               .mgr__std__lane22_strm0_data          ( mgr__std__lane22_strm0_data       ),      
               .mgr__std__lane22_strm0_data_valid    ( mgr__std__lane22_strm0_data_valid ),      
               .std__mgr__lane22_strm1_ready         ( std__mgr__lane22_strm1_ready      ),      
               .mgr__std__lane22_strm1_cntl          ( mgr__std__lane22_strm1_cntl       ),      
               .mgr__std__lane22_strm1_data          ( mgr__std__lane22_strm1_data       ),      
               .mgr__std__lane22_strm1_data_valid    ( mgr__std__lane22_strm1_data_valid ),      
               // Lane 23                 
               .std__mgr__lane23_strm0_ready         ( std__mgr__lane23_strm0_ready      ),      
               .mgr__std__lane23_strm0_cntl          ( mgr__std__lane23_strm0_cntl       ),      
               .mgr__std__lane23_strm0_data          ( mgr__std__lane23_strm0_data       ),      
               .mgr__std__lane23_strm0_data_valid    ( mgr__std__lane23_strm0_data_valid ),      
               .std__mgr__lane23_strm1_ready         ( std__mgr__lane23_strm1_ready      ),      
               .mgr__std__lane23_strm1_cntl          ( mgr__std__lane23_strm1_cntl       ),      
               .mgr__std__lane23_strm1_data          ( mgr__std__lane23_strm1_data       ),      
               .mgr__std__lane23_strm1_data_valid    ( mgr__std__lane23_strm1_data_valid ),      
               // Lane 24                 
               .std__mgr__lane24_strm0_ready         ( std__mgr__lane24_strm0_ready      ),      
               .mgr__std__lane24_strm0_cntl          ( mgr__std__lane24_strm0_cntl       ),      
               .mgr__std__lane24_strm0_data          ( mgr__std__lane24_strm0_data       ),      
               .mgr__std__lane24_strm0_data_valid    ( mgr__std__lane24_strm0_data_valid ),      
               .std__mgr__lane24_strm1_ready         ( std__mgr__lane24_strm1_ready      ),      
               .mgr__std__lane24_strm1_cntl          ( mgr__std__lane24_strm1_cntl       ),      
               .mgr__std__lane24_strm1_data          ( mgr__std__lane24_strm1_data       ),      
               .mgr__std__lane24_strm1_data_valid    ( mgr__std__lane24_strm1_data_valid ),      
               // Lane 25                 
               .std__mgr__lane25_strm0_ready         ( std__mgr__lane25_strm0_ready      ),      
               .mgr__std__lane25_strm0_cntl          ( mgr__std__lane25_strm0_cntl       ),      
               .mgr__std__lane25_strm0_data          ( mgr__std__lane25_strm0_data       ),      
               .mgr__std__lane25_strm0_data_valid    ( mgr__std__lane25_strm0_data_valid ),      
               .std__mgr__lane25_strm1_ready         ( std__mgr__lane25_strm1_ready      ),      
               .mgr__std__lane25_strm1_cntl          ( mgr__std__lane25_strm1_cntl       ),      
               .mgr__std__lane25_strm1_data          ( mgr__std__lane25_strm1_data       ),      
               .mgr__std__lane25_strm1_data_valid    ( mgr__std__lane25_strm1_data_valid ),      
               // Lane 26                 
               .std__mgr__lane26_strm0_ready         ( std__mgr__lane26_strm0_ready      ),      
               .mgr__std__lane26_strm0_cntl          ( mgr__std__lane26_strm0_cntl       ),      
               .mgr__std__lane26_strm0_data          ( mgr__std__lane26_strm0_data       ),      
               .mgr__std__lane26_strm0_data_valid    ( mgr__std__lane26_strm0_data_valid ),      
               .std__mgr__lane26_strm1_ready         ( std__mgr__lane26_strm1_ready      ),      
               .mgr__std__lane26_strm1_cntl          ( mgr__std__lane26_strm1_cntl       ),      
               .mgr__std__lane26_strm1_data          ( mgr__std__lane26_strm1_data       ),      
               .mgr__std__lane26_strm1_data_valid    ( mgr__std__lane26_strm1_data_valid ),      
               // Lane 27                 
               .std__mgr__lane27_strm0_ready         ( std__mgr__lane27_strm0_ready      ),      
               .mgr__std__lane27_strm0_cntl          ( mgr__std__lane27_strm0_cntl       ),      
               .mgr__std__lane27_strm0_data          ( mgr__std__lane27_strm0_data       ),      
               .mgr__std__lane27_strm0_data_valid    ( mgr__std__lane27_strm0_data_valid ),      
               .std__mgr__lane27_strm1_ready         ( std__mgr__lane27_strm1_ready      ),      
               .mgr__std__lane27_strm1_cntl          ( mgr__std__lane27_strm1_cntl       ),      
               .mgr__std__lane27_strm1_data          ( mgr__std__lane27_strm1_data       ),      
               .mgr__std__lane27_strm1_data_valid    ( mgr__std__lane27_strm1_data_valid ),      
               // Lane 28                 
               .std__mgr__lane28_strm0_ready         ( std__mgr__lane28_strm0_ready      ),      
               .mgr__std__lane28_strm0_cntl          ( mgr__std__lane28_strm0_cntl       ),      
               .mgr__std__lane28_strm0_data          ( mgr__std__lane28_strm0_data       ),      
               .mgr__std__lane28_strm0_data_valid    ( mgr__std__lane28_strm0_data_valid ),      
               .std__mgr__lane28_strm1_ready         ( std__mgr__lane28_strm1_ready      ),      
               .mgr__std__lane28_strm1_cntl          ( mgr__std__lane28_strm1_cntl       ),      
               .mgr__std__lane28_strm1_data          ( mgr__std__lane28_strm1_data       ),      
               .mgr__std__lane28_strm1_data_valid    ( mgr__std__lane28_strm1_data_valid ),      
               // Lane 29                 
               .std__mgr__lane29_strm0_ready         ( std__mgr__lane29_strm0_ready      ),      
               .mgr__std__lane29_strm0_cntl          ( mgr__std__lane29_strm0_cntl       ),      
               .mgr__std__lane29_strm0_data          ( mgr__std__lane29_strm0_data       ),      
               .mgr__std__lane29_strm0_data_valid    ( mgr__std__lane29_strm0_data_valid ),      
               .std__mgr__lane29_strm1_ready         ( std__mgr__lane29_strm1_ready      ),      
               .mgr__std__lane29_strm1_cntl          ( mgr__std__lane29_strm1_cntl       ),      
               .mgr__std__lane29_strm1_data          ( mgr__std__lane29_strm1_data       ),      
               .mgr__std__lane29_strm1_data_valid    ( mgr__std__lane29_strm1_data_valid ),      
               // Lane 30                 
               .std__mgr__lane30_strm0_ready         ( std__mgr__lane30_strm0_ready      ),      
               .mgr__std__lane30_strm0_cntl          ( mgr__std__lane30_strm0_cntl       ),      
               .mgr__std__lane30_strm0_data          ( mgr__std__lane30_strm0_data       ),      
               .mgr__std__lane30_strm0_data_valid    ( mgr__std__lane30_strm0_data_valid ),      
               .std__mgr__lane30_strm1_ready         ( std__mgr__lane30_strm1_ready      ),      
               .mgr__std__lane30_strm1_cntl          ( mgr__std__lane30_strm1_cntl       ),      
               .mgr__std__lane30_strm1_data          ( mgr__std__lane30_strm1_data       ),      
               .mgr__std__lane30_strm1_data_valid    ( mgr__std__lane30_strm1_data_valid ),      
               // Lane 31                 
               .std__mgr__lane31_strm0_ready         ( std__mgr__lane31_strm0_ready      ),      
               .mgr__std__lane31_strm0_cntl          ( mgr__std__lane31_strm0_cntl       ),      
               .mgr__std__lane31_strm0_data          ( mgr__std__lane31_strm0_data       ),      
               .mgr__std__lane31_strm0_data_valid    ( mgr__std__lane31_strm0_data_valid ),      
               .std__mgr__lane31_strm1_ready         ( std__mgr__lane31_strm1_ready      ),      
               .mgr__std__lane31_strm1_cntl          ( mgr__std__lane31_strm1_cntl       ),      
               .mgr__std__lane31_strm1_data          ( mgr__std__lane31_strm1_data       ),      
               .mgr__std__lane31_strm1_data_valid    ( mgr__std__lane31_strm1_data_valid ),      