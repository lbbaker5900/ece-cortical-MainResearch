
  // DMA accesses
        wire read_pause0        ;
        wire read_request0      ;
        wire read_access0       ;
        wire write_request0     ;
        wire write_access0      ;
        wire read_ready_strm0   ;  // ignore all requests until we deassert ready
        wire write_ready_strm0  ;  // ignore all requests until we deassert ready
        wire read_pause1        ;
        wire read_request1      ;
        wire read_access1       ;
        wire write_request1     ;
        wire write_access1      ;
        wire read_ready_strm1   ;  // ignore all requests until we deassert ready
        wire write_ready_strm1  ;  // ignore all requests until we deassert ready
        wire read_pause2        ;
        wire read_request2      ;
        wire read_access2       ;
        wire write_request2     ;
        wire write_access2      ;
        wire read_ready_strm2   ;  // ignore all requests until we deassert ready
        wire write_ready_strm2  ;  // ignore all requests until we deassert ready
        wire read_pause3        ;
        wire read_request3      ;
        wire read_access3       ;
        wire write_request3     ;
        wire write_access3      ;
        wire read_ready_strm3   ;  // ignore all requests until we deassert ready
        wire write_ready_strm3  ;  // ignore all requests until we deassert ready
        wire read_pause4        ;
        wire read_request4      ;
        wire read_access4       ;
        wire write_request4     ;
        wire write_access4      ;
        wire read_ready_strm4   ;  // ignore all requests until we deassert ready
        wire write_ready_strm4  ;  // ignore all requests until we deassert ready
        wire read_pause5        ;
        wire read_request5      ;
        wire read_access5       ;
        wire write_request5     ;
        wire write_access5      ;
        wire read_ready_strm5   ;  // ignore all requests until we deassert ready
        wire write_ready_strm5  ;  // ignore all requests until we deassert ready
        wire read_pause6        ;
        wire read_request6      ;
        wire read_access6       ;
        wire write_request6     ;
        wire write_access6      ;
        wire read_ready_strm6   ;  // ignore all requests until we deassert ready
        wire write_ready_strm6  ;  // ignore all requests until we deassert ready
        wire read_pause7        ;
        wire read_request7      ;
        wire read_access7       ;
        wire write_request7     ;
        wire write_access7      ;
        wire read_ready_strm7   ;  // ignore all requests until we deassert ready
        wire write_ready_strm7  ;  // ignore all requests until we deassert ready
        wire read_pause8        ;
        wire read_request8      ;
        wire read_access8       ;
        wire write_request8     ;
        wire write_access8      ;
        wire read_ready_strm8   ;  // ignore all requests until we deassert ready
        wire write_ready_strm8  ;  // ignore all requests until we deassert ready
        wire read_pause9        ;
        wire read_request9      ;
        wire read_access9       ;
        wire write_request9     ;
        wire write_access9      ;
        wire read_ready_strm9   ;  // ignore all requests until we deassert ready
        wire write_ready_strm9  ;  // ignore all requests until we deassert ready
        wire read_pause10        ;
        wire read_request10      ;
        wire read_access10       ;
        wire write_request10     ;
        wire write_access10      ;
        wire read_ready_strm10   ;  // ignore all requests until we deassert ready
        wire write_ready_strm10  ;  // ignore all requests until we deassert ready
        wire read_pause11        ;
        wire read_request11      ;
        wire read_access11       ;
        wire write_request11     ;
        wire write_access11      ;
        wire read_ready_strm11   ;  // ignore all requests until we deassert ready
        wire write_ready_strm11  ;  // ignore all requests until we deassert ready
        wire read_pause12        ;
        wire read_request12      ;
        wire read_access12       ;
        wire write_request12     ;
        wire write_access12      ;
        wire read_ready_strm12   ;  // ignore all requests until we deassert ready
        wire write_ready_strm12  ;  // ignore all requests until we deassert ready
        wire read_pause13        ;
        wire read_request13      ;
        wire read_access13       ;
        wire write_request13     ;
        wire write_access13      ;
        wire read_ready_strm13   ;  // ignore all requests until we deassert ready
        wire write_ready_strm13  ;  // ignore all requests until we deassert ready
        wire read_pause14        ;
        wire read_request14      ;
        wire read_access14       ;
        wire write_request14     ;
        wire write_access14      ;
        wire read_ready_strm14   ;  // ignore all requests until we deassert ready
        wire write_ready_strm14  ;  // ignore all requests until we deassert ready
        wire read_pause15        ;
        wire read_request15      ;
        wire read_access15       ;
        wire write_request15     ;
        wire write_access15      ;
        wire read_ready_strm15   ;  // ignore all requests until we deassert ready
        wire write_ready_strm15  ;  // ignore all requests until we deassert ready
        wire read_pause16        ;
        wire read_request16      ;
        wire read_access16       ;
        wire write_request16     ;
        wire write_access16      ;
        wire read_ready_strm16   ;  // ignore all requests until we deassert ready
        wire write_ready_strm16  ;  // ignore all requests until we deassert ready
        wire read_pause17        ;
        wire read_request17      ;
        wire read_access17       ;
        wire write_request17     ;
        wire write_access17      ;
        wire read_ready_strm17   ;  // ignore all requests until we deassert ready
        wire write_ready_strm17  ;  // ignore all requests until we deassert ready
        wire read_pause18        ;
        wire read_request18      ;
        wire read_access18       ;
        wire write_request18     ;
        wire write_access18      ;
        wire read_ready_strm18   ;  // ignore all requests until we deassert ready
        wire write_ready_strm18  ;  // ignore all requests until we deassert ready
        wire read_pause19        ;
        wire read_request19      ;
        wire read_access19       ;
        wire write_request19     ;
        wire write_access19      ;
        wire read_ready_strm19   ;  // ignore all requests until we deassert ready
        wire write_ready_strm19  ;  // ignore all requests until we deassert ready
        wire read_pause20        ;
        wire read_request20      ;
        wire read_access20       ;
        wire write_request20     ;
        wire write_access20      ;
        wire read_ready_strm20   ;  // ignore all requests until we deassert ready
        wire write_ready_strm20  ;  // ignore all requests until we deassert ready
        wire read_pause21        ;
        wire read_request21      ;
        wire read_access21       ;
        wire write_request21     ;
        wire write_access21      ;
        wire read_ready_strm21   ;  // ignore all requests until we deassert ready
        wire write_ready_strm21  ;  // ignore all requests until we deassert ready
        wire read_pause22        ;
        wire read_request22      ;
        wire read_access22       ;
        wire write_request22     ;
        wire write_access22      ;
        wire read_ready_strm22   ;  // ignore all requests until we deassert ready
        wire write_ready_strm22  ;  // ignore all requests until we deassert ready
        wire read_pause23        ;
        wire read_request23      ;
        wire read_access23       ;
        wire write_request23     ;
        wire write_access23      ;
        wire read_ready_strm23   ;  // ignore all requests until we deassert ready
        wire write_ready_strm23  ;  // ignore all requests until we deassert ready
        wire read_pause24        ;
        wire read_request24      ;
        wire read_access24       ;
        wire write_request24     ;
        wire write_access24      ;
        wire read_ready_strm24   ;  // ignore all requests until we deassert ready
        wire write_ready_strm24  ;  // ignore all requests until we deassert ready
        wire read_pause25        ;
        wire read_request25      ;
        wire read_access25       ;
        wire write_request25     ;
        wire write_access25      ;
        wire read_ready_strm25   ;  // ignore all requests until we deassert ready
        wire write_ready_strm25  ;  // ignore all requests until we deassert ready
        wire read_pause26        ;
        wire read_request26      ;
        wire read_access26       ;
        wire write_request26     ;
        wire write_access26      ;
        wire read_ready_strm26   ;  // ignore all requests until we deassert ready
        wire write_ready_strm26  ;  // ignore all requests until we deassert ready
        wire read_pause27        ;
        wire read_request27      ;
        wire read_access27       ;
        wire write_request27     ;
        wire write_access27      ;
        wire read_ready_strm27   ;  // ignore all requests until we deassert ready
        wire write_ready_strm27  ;  // ignore all requests until we deassert ready
        wire read_pause28        ;
        wire read_request28      ;
        wire read_access28       ;
        wire write_request28     ;
        wire write_access28      ;
        wire read_ready_strm28   ;  // ignore all requests until we deassert ready
        wire write_ready_strm28  ;  // ignore all requests until we deassert ready
        wire read_pause29        ;
        wire read_request29      ;
        wire read_access29       ;
        wire write_request29     ;
        wire write_access29      ;
        wire read_ready_strm29   ;  // ignore all requests until we deassert ready
        wire write_ready_strm29  ;  // ignore all requests until we deassert ready
        wire read_pause30        ;
        wire read_request30      ;
        wire read_access30       ;
        wire write_request30     ;
        wire write_access30      ;
        wire read_ready_strm30   ;  // ignore all requests until we deassert ready
        wire write_ready_strm30  ;  // ignore all requests until we deassert ready
        wire read_pause31        ;
        wire read_request31      ;
        wire read_access31       ;
        wire write_request31     ;
        wire write_access31      ;
        wire read_ready_strm31   ;  // ignore all requests until we deassert ready
        wire write_ready_strm31  ;  // ignore all requests until we deassert ready