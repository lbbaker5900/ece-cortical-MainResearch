
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__stu__valid        ( PeArray2Sys[0].pe__stu__valid             ),      
        .pe0__stu__cntl         ( PeArray2Sys[0].pe__stu__cntl              ),      
        .stu__pe0__ready        ( 1'b1     ),      
        //.stu__pe0__ready        ( PeArray2Sys[0].cb_test.stu__pe__ready     ),      
        .pe0__stu__type         ( PeArray2Sys[0].pe__stu__type              ),      
        .pe0__stu__data         ( PeArray2Sys[0].pe__stu__data              ),      
        .pe0__stu__oob_data     ( PeArray2Sys[0].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__stu__valid        ( PeArray2Sys[1].pe__stu__valid             ),      
        .pe1__stu__cntl         ( PeArray2Sys[1].pe__stu__cntl              ),      
        .stu__pe1__ready        ( 1'b1     ),      
        //.stu__pe1__ready        ( PeArray2Sys[1].cb_test.stu__pe__ready     ),      
        .pe1__stu__type         ( PeArray2Sys[1].pe__stu__type              ),      
        .pe1__stu__data         ( PeArray2Sys[1].pe__stu__data              ),      
        .pe1__stu__oob_data     ( PeArray2Sys[1].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__stu__valid        ( PeArray2Sys[2].pe__stu__valid             ),      
        .pe2__stu__cntl         ( PeArray2Sys[2].pe__stu__cntl              ),      
        .stu__pe2__ready        ( 1'b1     ),      
        //.stu__pe2__ready        ( PeArray2Sys[2].cb_test.stu__pe__ready     ),      
        .pe2__stu__type         ( PeArray2Sys[2].pe__stu__type              ),      
        .pe2__stu__data         ( PeArray2Sys[2].pe__stu__data              ),      
        .pe2__stu__oob_data     ( PeArray2Sys[2].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__stu__valid        ( PeArray2Sys[3].pe__stu__valid             ),      
        .pe3__stu__cntl         ( PeArray2Sys[3].pe__stu__cntl              ),      
        .stu__pe3__ready        ( 1'b1     ),      
        //.stu__pe3__ready        ( PeArray2Sys[3].cb_test.stu__pe__ready     ),      
        .pe3__stu__type         ( PeArray2Sys[3].pe__stu__type              ),      
        .pe3__stu__data         ( PeArray2Sys[3].pe__stu__data              ),      
        .pe3__stu__oob_data     ( PeArray2Sys[3].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__stu__valid        ( PeArray2Sys[4].pe__stu__valid             ),      
        .pe4__stu__cntl         ( PeArray2Sys[4].pe__stu__cntl              ),      
        .stu__pe4__ready        ( 1'b1     ),      
        //.stu__pe4__ready        ( PeArray2Sys[4].cb_test.stu__pe__ready     ),      
        .pe4__stu__type         ( PeArray2Sys[4].pe__stu__type              ),      
        .pe4__stu__data         ( PeArray2Sys[4].pe__stu__data              ),      
        .pe4__stu__oob_data     ( PeArray2Sys[4].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__stu__valid        ( PeArray2Sys[5].pe__stu__valid             ),      
        .pe5__stu__cntl         ( PeArray2Sys[5].pe__stu__cntl              ),      
        .stu__pe5__ready        ( 1'b1     ),      
        //.stu__pe5__ready        ( PeArray2Sys[5].cb_test.stu__pe__ready     ),      
        .pe5__stu__type         ( PeArray2Sys[5].pe__stu__type              ),      
        .pe5__stu__data         ( PeArray2Sys[5].pe__stu__data              ),      
        .pe5__stu__oob_data     ( PeArray2Sys[5].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__stu__valid        ( PeArray2Sys[6].pe__stu__valid             ),      
        .pe6__stu__cntl         ( PeArray2Sys[6].pe__stu__cntl              ),      
        .stu__pe6__ready        ( 1'b1     ),      
        //.stu__pe6__ready        ( PeArray2Sys[6].cb_test.stu__pe__ready     ),      
        .pe6__stu__type         ( PeArray2Sys[6].pe__stu__type              ),      
        .pe6__stu__data         ( PeArray2Sys[6].pe__stu__data              ),      
        .pe6__stu__oob_data     ( PeArray2Sys[6].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__stu__valid        ( PeArray2Sys[7].pe__stu__valid             ),      
        .pe7__stu__cntl         ( PeArray2Sys[7].pe__stu__cntl              ),      
        .stu__pe7__ready        ( 1'b1     ),      
        //.stu__pe7__ready        ( PeArray2Sys[7].cb_test.stu__pe__ready     ),      
        .pe7__stu__type         ( PeArray2Sys[7].pe__stu__type              ),      
        .pe7__stu__data         ( PeArray2Sys[7].pe__stu__data              ),      
        .pe7__stu__oob_data     ( PeArray2Sys[7].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__stu__valid        ( PeArray2Sys[8].pe__stu__valid             ),      
        .pe8__stu__cntl         ( PeArray2Sys[8].pe__stu__cntl              ),      
        .stu__pe8__ready        ( 1'b1     ),      
        //.stu__pe8__ready        ( PeArray2Sys[8].cb_test.stu__pe__ready     ),      
        .pe8__stu__type         ( PeArray2Sys[8].pe__stu__type              ),      
        .pe8__stu__data         ( PeArray2Sys[8].pe__stu__data              ),      
        .pe8__stu__oob_data     ( PeArray2Sys[8].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__stu__valid        ( PeArray2Sys[9].pe__stu__valid             ),      
        .pe9__stu__cntl         ( PeArray2Sys[9].pe__stu__cntl              ),      
        .stu__pe9__ready        ( 1'b1     ),      
        //.stu__pe9__ready        ( PeArray2Sys[9].cb_test.stu__pe__ready     ),      
        .pe9__stu__type         ( PeArray2Sys[9].pe__stu__type              ),      
        .pe9__stu__data         ( PeArray2Sys[9].pe__stu__data              ),      
        .pe9__stu__oob_data     ( PeArray2Sys[9].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__stu__valid        ( PeArray2Sys[10].pe__stu__valid             ),      
        .pe10__stu__cntl         ( PeArray2Sys[10].pe__stu__cntl              ),      
        .stu__pe10__ready        ( 1'b1     ),      
        //.stu__pe10__ready        ( PeArray2Sys[10].cb_test.stu__pe__ready     ),      
        .pe10__stu__type         ( PeArray2Sys[10].pe__stu__type              ),      
        .pe10__stu__data         ( PeArray2Sys[10].pe__stu__data              ),      
        .pe10__stu__oob_data     ( PeArray2Sys[10].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__stu__valid        ( PeArray2Sys[11].pe__stu__valid             ),      
        .pe11__stu__cntl         ( PeArray2Sys[11].pe__stu__cntl              ),      
        .stu__pe11__ready        ( 1'b1     ),      
        //.stu__pe11__ready        ( PeArray2Sys[11].cb_test.stu__pe__ready     ),      
        .pe11__stu__type         ( PeArray2Sys[11].pe__stu__type              ),      
        .pe11__stu__data         ( PeArray2Sys[11].pe__stu__data              ),      
        .pe11__stu__oob_data     ( PeArray2Sys[11].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__stu__valid        ( PeArray2Sys[12].pe__stu__valid             ),      
        .pe12__stu__cntl         ( PeArray2Sys[12].pe__stu__cntl              ),      
        .stu__pe12__ready        ( 1'b1     ),      
        //.stu__pe12__ready        ( PeArray2Sys[12].cb_test.stu__pe__ready     ),      
        .pe12__stu__type         ( PeArray2Sys[12].pe__stu__type              ),      
        .pe12__stu__data         ( PeArray2Sys[12].pe__stu__data              ),      
        .pe12__stu__oob_data     ( PeArray2Sys[12].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__stu__valid        ( PeArray2Sys[13].pe__stu__valid             ),      
        .pe13__stu__cntl         ( PeArray2Sys[13].pe__stu__cntl              ),      
        .stu__pe13__ready        ( 1'b1     ),      
        //.stu__pe13__ready        ( PeArray2Sys[13].cb_test.stu__pe__ready     ),      
        .pe13__stu__type         ( PeArray2Sys[13].pe__stu__type              ),      
        .pe13__stu__data         ( PeArray2Sys[13].pe__stu__data              ),      
        .pe13__stu__oob_data     ( PeArray2Sys[13].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__stu__valid        ( PeArray2Sys[14].pe__stu__valid             ),      
        .pe14__stu__cntl         ( PeArray2Sys[14].pe__stu__cntl              ),      
        .stu__pe14__ready        ( 1'b1     ),      
        //.stu__pe14__ready        ( PeArray2Sys[14].cb_test.stu__pe__ready     ),      
        .pe14__stu__type         ( PeArray2Sys[14].pe__stu__type              ),      
        .pe14__stu__data         ( PeArray2Sys[14].pe__stu__data              ),      
        .pe14__stu__oob_data     ( PeArray2Sys[14].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__stu__valid        ( PeArray2Sys[15].pe__stu__valid             ),      
        .pe15__stu__cntl         ( PeArray2Sys[15].pe__stu__cntl              ),      
        .stu__pe15__ready        ( 1'b1     ),      
        //.stu__pe15__ready        ( PeArray2Sys[15].cb_test.stu__pe__ready     ),      
        .pe15__stu__type         ( PeArray2Sys[15].pe__stu__type              ),      
        .pe15__stu__data         ( PeArray2Sys[15].pe__stu__data              ),      
        .pe15__stu__oob_data     ( PeArray2Sys[15].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__stu__valid        ( PeArray2Sys[16].pe__stu__valid             ),      
        .pe16__stu__cntl         ( PeArray2Sys[16].pe__stu__cntl              ),      
        .stu__pe16__ready        ( 1'b1     ),      
        //.stu__pe16__ready        ( PeArray2Sys[16].cb_test.stu__pe__ready     ),      
        .pe16__stu__type         ( PeArray2Sys[16].pe__stu__type              ),      
        .pe16__stu__data         ( PeArray2Sys[16].pe__stu__data              ),      
        .pe16__stu__oob_data     ( PeArray2Sys[16].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__stu__valid        ( PeArray2Sys[17].pe__stu__valid             ),      
        .pe17__stu__cntl         ( PeArray2Sys[17].pe__stu__cntl              ),      
        .stu__pe17__ready        ( 1'b1     ),      
        //.stu__pe17__ready        ( PeArray2Sys[17].cb_test.stu__pe__ready     ),      
        .pe17__stu__type         ( PeArray2Sys[17].pe__stu__type              ),      
        .pe17__stu__data         ( PeArray2Sys[17].pe__stu__data              ),      
        .pe17__stu__oob_data     ( PeArray2Sys[17].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__stu__valid        ( PeArray2Sys[18].pe__stu__valid             ),      
        .pe18__stu__cntl         ( PeArray2Sys[18].pe__stu__cntl              ),      
        .stu__pe18__ready        ( 1'b1     ),      
        //.stu__pe18__ready        ( PeArray2Sys[18].cb_test.stu__pe__ready     ),      
        .pe18__stu__type         ( PeArray2Sys[18].pe__stu__type              ),      
        .pe18__stu__data         ( PeArray2Sys[18].pe__stu__data              ),      
        .pe18__stu__oob_data     ( PeArray2Sys[18].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__stu__valid        ( PeArray2Sys[19].pe__stu__valid             ),      
        .pe19__stu__cntl         ( PeArray2Sys[19].pe__stu__cntl              ),      
        .stu__pe19__ready        ( 1'b1     ),      
        //.stu__pe19__ready        ( PeArray2Sys[19].cb_test.stu__pe__ready     ),      
        .pe19__stu__type         ( PeArray2Sys[19].pe__stu__type              ),      
        .pe19__stu__data         ( PeArray2Sys[19].pe__stu__data              ),      
        .pe19__stu__oob_data     ( PeArray2Sys[19].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__stu__valid        ( PeArray2Sys[20].pe__stu__valid             ),      
        .pe20__stu__cntl         ( PeArray2Sys[20].pe__stu__cntl              ),      
        .stu__pe20__ready        ( 1'b1     ),      
        //.stu__pe20__ready        ( PeArray2Sys[20].cb_test.stu__pe__ready     ),      
        .pe20__stu__type         ( PeArray2Sys[20].pe__stu__type              ),      
        .pe20__stu__data         ( PeArray2Sys[20].pe__stu__data              ),      
        .pe20__stu__oob_data     ( PeArray2Sys[20].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__stu__valid        ( PeArray2Sys[21].pe__stu__valid             ),      
        .pe21__stu__cntl         ( PeArray2Sys[21].pe__stu__cntl              ),      
        .stu__pe21__ready        ( 1'b1     ),      
        //.stu__pe21__ready        ( PeArray2Sys[21].cb_test.stu__pe__ready     ),      
        .pe21__stu__type         ( PeArray2Sys[21].pe__stu__type              ),      
        .pe21__stu__data         ( PeArray2Sys[21].pe__stu__data              ),      
        .pe21__stu__oob_data     ( PeArray2Sys[21].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__stu__valid        ( PeArray2Sys[22].pe__stu__valid             ),      
        .pe22__stu__cntl         ( PeArray2Sys[22].pe__stu__cntl              ),      
        .stu__pe22__ready        ( 1'b1     ),      
        //.stu__pe22__ready        ( PeArray2Sys[22].cb_test.stu__pe__ready     ),      
        .pe22__stu__type         ( PeArray2Sys[22].pe__stu__type              ),      
        .pe22__stu__data         ( PeArray2Sys[22].pe__stu__data              ),      
        .pe22__stu__oob_data     ( PeArray2Sys[22].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__stu__valid        ( PeArray2Sys[23].pe__stu__valid             ),      
        .pe23__stu__cntl         ( PeArray2Sys[23].pe__stu__cntl              ),      
        .stu__pe23__ready        ( 1'b1     ),      
        //.stu__pe23__ready        ( PeArray2Sys[23].cb_test.stu__pe__ready     ),      
        .pe23__stu__type         ( PeArray2Sys[23].pe__stu__type              ),      
        .pe23__stu__data         ( PeArray2Sys[23].pe__stu__data              ),      
        .pe23__stu__oob_data     ( PeArray2Sys[23].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__stu__valid        ( PeArray2Sys[24].pe__stu__valid             ),      
        .pe24__stu__cntl         ( PeArray2Sys[24].pe__stu__cntl              ),      
        .stu__pe24__ready        ( 1'b1     ),      
        //.stu__pe24__ready        ( PeArray2Sys[24].cb_test.stu__pe__ready     ),      
        .pe24__stu__type         ( PeArray2Sys[24].pe__stu__type              ),      
        .pe24__stu__data         ( PeArray2Sys[24].pe__stu__data              ),      
        .pe24__stu__oob_data     ( PeArray2Sys[24].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__stu__valid        ( PeArray2Sys[25].pe__stu__valid             ),      
        .pe25__stu__cntl         ( PeArray2Sys[25].pe__stu__cntl              ),      
        .stu__pe25__ready        ( 1'b1     ),      
        //.stu__pe25__ready        ( PeArray2Sys[25].cb_test.stu__pe__ready     ),      
        .pe25__stu__type         ( PeArray2Sys[25].pe__stu__type              ),      
        .pe25__stu__data         ( PeArray2Sys[25].pe__stu__data              ),      
        .pe25__stu__oob_data     ( PeArray2Sys[25].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__stu__valid        ( PeArray2Sys[26].pe__stu__valid             ),      
        .pe26__stu__cntl         ( PeArray2Sys[26].pe__stu__cntl              ),      
        .stu__pe26__ready        ( 1'b1     ),      
        //.stu__pe26__ready        ( PeArray2Sys[26].cb_test.stu__pe__ready     ),      
        .pe26__stu__type         ( PeArray2Sys[26].pe__stu__type              ),      
        .pe26__stu__data         ( PeArray2Sys[26].pe__stu__data              ),      
        .pe26__stu__oob_data     ( PeArray2Sys[26].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__stu__valid        ( PeArray2Sys[27].pe__stu__valid             ),      
        .pe27__stu__cntl         ( PeArray2Sys[27].pe__stu__cntl              ),      
        .stu__pe27__ready        ( 1'b1     ),      
        //.stu__pe27__ready        ( PeArray2Sys[27].cb_test.stu__pe__ready     ),      
        .pe27__stu__type         ( PeArray2Sys[27].pe__stu__type              ),      
        .pe27__stu__data         ( PeArray2Sys[27].pe__stu__data              ),      
        .pe27__stu__oob_data     ( PeArray2Sys[27].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__stu__valid        ( PeArray2Sys[28].pe__stu__valid             ),      
        .pe28__stu__cntl         ( PeArray2Sys[28].pe__stu__cntl              ),      
        .stu__pe28__ready        ( 1'b1     ),      
        //.stu__pe28__ready        ( PeArray2Sys[28].cb_test.stu__pe__ready     ),      
        .pe28__stu__type         ( PeArray2Sys[28].pe__stu__type              ),      
        .pe28__stu__data         ( PeArray2Sys[28].pe__stu__data              ),      
        .pe28__stu__oob_data     ( PeArray2Sys[28].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__stu__valid        ( PeArray2Sys[29].pe__stu__valid             ),      
        .pe29__stu__cntl         ( PeArray2Sys[29].pe__stu__cntl              ),      
        .stu__pe29__ready        ( 1'b1     ),      
        //.stu__pe29__ready        ( PeArray2Sys[29].cb_test.stu__pe__ready     ),      
        .pe29__stu__type         ( PeArray2Sys[29].pe__stu__type              ),      
        .pe29__stu__data         ( PeArray2Sys[29].pe__stu__data              ),      
        .pe29__stu__oob_data     ( PeArray2Sys[29].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__stu__valid        ( PeArray2Sys[30].pe__stu__valid             ),      
        .pe30__stu__cntl         ( PeArray2Sys[30].pe__stu__cntl              ),      
        .stu__pe30__ready        ( 1'b1     ),      
        //.stu__pe30__ready        ( PeArray2Sys[30].cb_test.stu__pe__ready     ),      
        .pe30__stu__type         ( PeArray2Sys[30].pe__stu__type              ),      
        .pe30__stu__data         ( PeArray2Sys[30].pe__stu__data              ),      
        .pe30__stu__oob_data     ( PeArray2Sys[30].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__stu__valid        ( PeArray2Sys[31].pe__stu__valid             ),      
        .pe31__stu__cntl         ( PeArray2Sys[31].pe__stu__cntl              ),      
        .stu__pe31__ready        ( 1'b1     ),      
        //.stu__pe31__ready        ( PeArray2Sys[31].cb_test.stu__pe__ready     ),      
        .pe31__stu__type         ( PeArray2Sys[31].pe__stu__type              ),      
        .pe31__stu__data         ( PeArray2Sys[31].pe__stu__data              ),      
        .pe31__stu__oob_data     ( PeArray2Sys[31].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__stu__valid        ( PeArray2Sys[32].pe__stu__valid             ),      
        .pe32__stu__cntl         ( PeArray2Sys[32].pe__stu__cntl              ),      
        .stu__pe32__ready        ( 1'b1     ),      
        //.stu__pe32__ready        ( PeArray2Sys[32].cb_test.stu__pe__ready     ),      
        .pe32__stu__type         ( PeArray2Sys[32].pe__stu__type              ),      
        .pe32__stu__data         ( PeArray2Sys[32].pe__stu__data              ),      
        .pe32__stu__oob_data     ( PeArray2Sys[32].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__stu__valid        ( PeArray2Sys[33].pe__stu__valid             ),      
        .pe33__stu__cntl         ( PeArray2Sys[33].pe__stu__cntl              ),      
        .stu__pe33__ready        ( 1'b1     ),      
        //.stu__pe33__ready        ( PeArray2Sys[33].cb_test.stu__pe__ready     ),      
        .pe33__stu__type         ( PeArray2Sys[33].pe__stu__type              ),      
        .pe33__stu__data         ( PeArray2Sys[33].pe__stu__data              ),      
        .pe33__stu__oob_data     ( PeArray2Sys[33].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__stu__valid        ( PeArray2Sys[34].pe__stu__valid             ),      
        .pe34__stu__cntl         ( PeArray2Sys[34].pe__stu__cntl              ),      
        .stu__pe34__ready        ( 1'b1     ),      
        //.stu__pe34__ready        ( PeArray2Sys[34].cb_test.stu__pe__ready     ),      
        .pe34__stu__type         ( PeArray2Sys[34].pe__stu__type              ),      
        .pe34__stu__data         ( PeArray2Sys[34].pe__stu__data              ),      
        .pe34__stu__oob_data     ( PeArray2Sys[34].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__stu__valid        ( PeArray2Sys[35].pe__stu__valid             ),      
        .pe35__stu__cntl         ( PeArray2Sys[35].pe__stu__cntl              ),      
        .stu__pe35__ready        ( 1'b1     ),      
        //.stu__pe35__ready        ( PeArray2Sys[35].cb_test.stu__pe__ready     ),      
        .pe35__stu__type         ( PeArray2Sys[35].pe__stu__type              ),      
        .pe35__stu__data         ( PeArray2Sys[35].pe__stu__data              ),      
        .pe35__stu__oob_data     ( PeArray2Sys[35].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__stu__valid        ( PeArray2Sys[36].pe__stu__valid             ),      
        .pe36__stu__cntl         ( PeArray2Sys[36].pe__stu__cntl              ),      
        .stu__pe36__ready        ( 1'b1     ),      
        //.stu__pe36__ready        ( PeArray2Sys[36].cb_test.stu__pe__ready     ),      
        .pe36__stu__type         ( PeArray2Sys[36].pe__stu__type              ),      
        .pe36__stu__data         ( PeArray2Sys[36].pe__stu__data              ),      
        .pe36__stu__oob_data     ( PeArray2Sys[36].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__stu__valid        ( PeArray2Sys[37].pe__stu__valid             ),      
        .pe37__stu__cntl         ( PeArray2Sys[37].pe__stu__cntl              ),      
        .stu__pe37__ready        ( 1'b1     ),      
        //.stu__pe37__ready        ( PeArray2Sys[37].cb_test.stu__pe__ready     ),      
        .pe37__stu__type         ( PeArray2Sys[37].pe__stu__type              ),      
        .pe37__stu__data         ( PeArray2Sys[37].pe__stu__data              ),      
        .pe37__stu__oob_data     ( PeArray2Sys[37].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__stu__valid        ( PeArray2Sys[38].pe__stu__valid             ),      
        .pe38__stu__cntl         ( PeArray2Sys[38].pe__stu__cntl              ),      
        .stu__pe38__ready        ( 1'b1     ),      
        //.stu__pe38__ready        ( PeArray2Sys[38].cb_test.stu__pe__ready     ),      
        .pe38__stu__type         ( PeArray2Sys[38].pe__stu__type              ),      
        .pe38__stu__data         ( PeArray2Sys[38].pe__stu__data              ),      
        .pe38__stu__oob_data     ( PeArray2Sys[38].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__stu__valid        ( PeArray2Sys[39].pe__stu__valid             ),      
        .pe39__stu__cntl         ( PeArray2Sys[39].pe__stu__cntl              ),      
        .stu__pe39__ready        ( 1'b1     ),      
        //.stu__pe39__ready        ( PeArray2Sys[39].cb_test.stu__pe__ready     ),      
        .pe39__stu__type         ( PeArray2Sys[39].pe__stu__type              ),      
        .pe39__stu__data         ( PeArray2Sys[39].pe__stu__data              ),      
        .pe39__stu__oob_data     ( PeArray2Sys[39].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__stu__valid        ( PeArray2Sys[40].pe__stu__valid             ),      
        .pe40__stu__cntl         ( PeArray2Sys[40].pe__stu__cntl              ),      
        .stu__pe40__ready        ( 1'b1     ),      
        //.stu__pe40__ready        ( PeArray2Sys[40].cb_test.stu__pe__ready     ),      
        .pe40__stu__type         ( PeArray2Sys[40].pe__stu__type              ),      
        .pe40__stu__data         ( PeArray2Sys[40].pe__stu__data              ),      
        .pe40__stu__oob_data     ( PeArray2Sys[40].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__stu__valid        ( PeArray2Sys[41].pe__stu__valid             ),      
        .pe41__stu__cntl         ( PeArray2Sys[41].pe__stu__cntl              ),      
        .stu__pe41__ready        ( 1'b1     ),      
        //.stu__pe41__ready        ( PeArray2Sys[41].cb_test.stu__pe__ready     ),      
        .pe41__stu__type         ( PeArray2Sys[41].pe__stu__type              ),      
        .pe41__stu__data         ( PeArray2Sys[41].pe__stu__data              ),      
        .pe41__stu__oob_data     ( PeArray2Sys[41].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__stu__valid        ( PeArray2Sys[42].pe__stu__valid             ),      
        .pe42__stu__cntl         ( PeArray2Sys[42].pe__stu__cntl              ),      
        .stu__pe42__ready        ( 1'b1     ),      
        //.stu__pe42__ready        ( PeArray2Sys[42].cb_test.stu__pe__ready     ),      
        .pe42__stu__type         ( PeArray2Sys[42].pe__stu__type              ),      
        .pe42__stu__data         ( PeArray2Sys[42].pe__stu__data              ),      
        .pe42__stu__oob_data     ( PeArray2Sys[42].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__stu__valid        ( PeArray2Sys[43].pe__stu__valid             ),      
        .pe43__stu__cntl         ( PeArray2Sys[43].pe__stu__cntl              ),      
        .stu__pe43__ready        ( 1'b1     ),      
        //.stu__pe43__ready        ( PeArray2Sys[43].cb_test.stu__pe__ready     ),      
        .pe43__stu__type         ( PeArray2Sys[43].pe__stu__type              ),      
        .pe43__stu__data         ( PeArray2Sys[43].pe__stu__data              ),      
        .pe43__stu__oob_data     ( PeArray2Sys[43].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__stu__valid        ( PeArray2Sys[44].pe__stu__valid             ),      
        .pe44__stu__cntl         ( PeArray2Sys[44].pe__stu__cntl              ),      
        .stu__pe44__ready        ( 1'b1     ),      
        //.stu__pe44__ready        ( PeArray2Sys[44].cb_test.stu__pe__ready     ),      
        .pe44__stu__type         ( PeArray2Sys[44].pe__stu__type              ),      
        .pe44__stu__data         ( PeArray2Sys[44].pe__stu__data              ),      
        .pe44__stu__oob_data     ( PeArray2Sys[44].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__stu__valid        ( PeArray2Sys[45].pe__stu__valid             ),      
        .pe45__stu__cntl         ( PeArray2Sys[45].pe__stu__cntl              ),      
        .stu__pe45__ready        ( 1'b1     ),      
        //.stu__pe45__ready        ( PeArray2Sys[45].cb_test.stu__pe__ready     ),      
        .pe45__stu__type         ( PeArray2Sys[45].pe__stu__type              ),      
        .pe45__stu__data         ( PeArray2Sys[45].pe__stu__data              ),      
        .pe45__stu__oob_data     ( PeArray2Sys[45].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__stu__valid        ( PeArray2Sys[46].pe__stu__valid             ),      
        .pe46__stu__cntl         ( PeArray2Sys[46].pe__stu__cntl              ),      
        .stu__pe46__ready        ( 1'b1     ),      
        //.stu__pe46__ready        ( PeArray2Sys[46].cb_test.stu__pe__ready     ),      
        .pe46__stu__type         ( PeArray2Sys[46].pe__stu__type              ),      
        .pe46__stu__data         ( PeArray2Sys[46].pe__stu__data              ),      
        .pe46__stu__oob_data     ( PeArray2Sys[46].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__stu__valid        ( PeArray2Sys[47].pe__stu__valid             ),      
        .pe47__stu__cntl         ( PeArray2Sys[47].pe__stu__cntl              ),      
        .stu__pe47__ready        ( 1'b1     ),      
        //.stu__pe47__ready        ( PeArray2Sys[47].cb_test.stu__pe__ready     ),      
        .pe47__stu__type         ( PeArray2Sys[47].pe__stu__type              ),      
        .pe47__stu__data         ( PeArray2Sys[47].pe__stu__data              ),      
        .pe47__stu__oob_data     ( PeArray2Sys[47].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__stu__valid        ( PeArray2Sys[48].pe__stu__valid             ),      
        .pe48__stu__cntl         ( PeArray2Sys[48].pe__stu__cntl              ),      
        .stu__pe48__ready        ( 1'b1     ),      
        //.stu__pe48__ready        ( PeArray2Sys[48].cb_test.stu__pe__ready     ),      
        .pe48__stu__type         ( PeArray2Sys[48].pe__stu__type              ),      
        .pe48__stu__data         ( PeArray2Sys[48].pe__stu__data              ),      
        .pe48__stu__oob_data     ( PeArray2Sys[48].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__stu__valid        ( PeArray2Sys[49].pe__stu__valid             ),      
        .pe49__stu__cntl         ( PeArray2Sys[49].pe__stu__cntl              ),      
        .stu__pe49__ready        ( 1'b1     ),      
        //.stu__pe49__ready        ( PeArray2Sys[49].cb_test.stu__pe__ready     ),      
        .pe49__stu__type         ( PeArray2Sys[49].pe__stu__type              ),      
        .pe49__stu__data         ( PeArray2Sys[49].pe__stu__data              ),      
        .pe49__stu__oob_data     ( PeArray2Sys[49].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__stu__valid        ( PeArray2Sys[50].pe__stu__valid             ),      
        .pe50__stu__cntl         ( PeArray2Sys[50].pe__stu__cntl              ),      
        .stu__pe50__ready        ( 1'b1     ),      
        //.stu__pe50__ready        ( PeArray2Sys[50].cb_test.stu__pe__ready     ),      
        .pe50__stu__type         ( PeArray2Sys[50].pe__stu__type              ),      
        .pe50__stu__data         ( PeArray2Sys[50].pe__stu__data              ),      
        .pe50__stu__oob_data     ( PeArray2Sys[50].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__stu__valid        ( PeArray2Sys[51].pe__stu__valid             ),      
        .pe51__stu__cntl         ( PeArray2Sys[51].pe__stu__cntl              ),      
        .stu__pe51__ready        ( 1'b1     ),      
        //.stu__pe51__ready        ( PeArray2Sys[51].cb_test.stu__pe__ready     ),      
        .pe51__stu__type         ( PeArray2Sys[51].pe__stu__type              ),      
        .pe51__stu__data         ( PeArray2Sys[51].pe__stu__data              ),      
        .pe51__stu__oob_data     ( PeArray2Sys[51].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__stu__valid        ( PeArray2Sys[52].pe__stu__valid             ),      
        .pe52__stu__cntl         ( PeArray2Sys[52].pe__stu__cntl              ),      
        .stu__pe52__ready        ( 1'b1     ),      
        //.stu__pe52__ready        ( PeArray2Sys[52].cb_test.stu__pe__ready     ),      
        .pe52__stu__type         ( PeArray2Sys[52].pe__stu__type              ),      
        .pe52__stu__data         ( PeArray2Sys[52].pe__stu__data              ),      
        .pe52__stu__oob_data     ( PeArray2Sys[52].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__stu__valid        ( PeArray2Sys[53].pe__stu__valid             ),      
        .pe53__stu__cntl         ( PeArray2Sys[53].pe__stu__cntl              ),      
        .stu__pe53__ready        ( 1'b1     ),      
        //.stu__pe53__ready        ( PeArray2Sys[53].cb_test.stu__pe__ready     ),      
        .pe53__stu__type         ( PeArray2Sys[53].pe__stu__type              ),      
        .pe53__stu__data         ( PeArray2Sys[53].pe__stu__data              ),      
        .pe53__stu__oob_data     ( PeArray2Sys[53].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__stu__valid        ( PeArray2Sys[54].pe__stu__valid             ),      
        .pe54__stu__cntl         ( PeArray2Sys[54].pe__stu__cntl              ),      
        .stu__pe54__ready        ( 1'b1     ),      
        //.stu__pe54__ready        ( PeArray2Sys[54].cb_test.stu__pe__ready     ),      
        .pe54__stu__type         ( PeArray2Sys[54].pe__stu__type              ),      
        .pe54__stu__data         ( PeArray2Sys[54].pe__stu__data              ),      
        .pe54__stu__oob_data     ( PeArray2Sys[54].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__stu__valid        ( PeArray2Sys[55].pe__stu__valid             ),      
        .pe55__stu__cntl         ( PeArray2Sys[55].pe__stu__cntl              ),      
        .stu__pe55__ready        ( 1'b1     ),      
        //.stu__pe55__ready        ( PeArray2Sys[55].cb_test.stu__pe__ready     ),      
        .pe55__stu__type         ( PeArray2Sys[55].pe__stu__type              ),      
        .pe55__stu__data         ( PeArray2Sys[55].pe__stu__data              ),      
        .pe55__stu__oob_data     ( PeArray2Sys[55].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__stu__valid        ( PeArray2Sys[56].pe__stu__valid             ),      
        .pe56__stu__cntl         ( PeArray2Sys[56].pe__stu__cntl              ),      
        .stu__pe56__ready        ( 1'b1     ),      
        //.stu__pe56__ready        ( PeArray2Sys[56].cb_test.stu__pe__ready     ),      
        .pe56__stu__type         ( PeArray2Sys[56].pe__stu__type              ),      
        .pe56__stu__data         ( PeArray2Sys[56].pe__stu__data              ),      
        .pe56__stu__oob_data     ( PeArray2Sys[56].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__stu__valid        ( PeArray2Sys[57].pe__stu__valid             ),      
        .pe57__stu__cntl         ( PeArray2Sys[57].pe__stu__cntl              ),      
        .stu__pe57__ready        ( 1'b1     ),      
        //.stu__pe57__ready        ( PeArray2Sys[57].cb_test.stu__pe__ready     ),      
        .pe57__stu__type         ( PeArray2Sys[57].pe__stu__type              ),      
        .pe57__stu__data         ( PeArray2Sys[57].pe__stu__data              ),      
        .pe57__stu__oob_data     ( PeArray2Sys[57].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__stu__valid        ( PeArray2Sys[58].pe__stu__valid             ),      
        .pe58__stu__cntl         ( PeArray2Sys[58].pe__stu__cntl              ),      
        .stu__pe58__ready        ( 1'b1     ),      
        //.stu__pe58__ready        ( PeArray2Sys[58].cb_test.stu__pe__ready     ),      
        .pe58__stu__type         ( PeArray2Sys[58].pe__stu__type              ),      
        .pe58__stu__data         ( PeArray2Sys[58].pe__stu__data              ),      
        .pe58__stu__oob_data     ( PeArray2Sys[58].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__stu__valid        ( PeArray2Sys[59].pe__stu__valid             ),      
        .pe59__stu__cntl         ( PeArray2Sys[59].pe__stu__cntl              ),      
        .stu__pe59__ready        ( 1'b1     ),      
        //.stu__pe59__ready        ( PeArray2Sys[59].cb_test.stu__pe__ready     ),      
        .pe59__stu__type         ( PeArray2Sys[59].pe__stu__type              ),      
        .pe59__stu__data         ( PeArray2Sys[59].pe__stu__data              ),      
        .pe59__stu__oob_data     ( PeArray2Sys[59].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__stu__valid        ( PeArray2Sys[60].pe__stu__valid             ),      
        .pe60__stu__cntl         ( PeArray2Sys[60].pe__stu__cntl              ),      
        .stu__pe60__ready        ( 1'b1     ),      
        //.stu__pe60__ready        ( PeArray2Sys[60].cb_test.stu__pe__ready     ),      
        .pe60__stu__type         ( PeArray2Sys[60].pe__stu__type              ),      
        .pe60__stu__data         ( PeArray2Sys[60].pe__stu__data              ),      
        .pe60__stu__oob_data     ( PeArray2Sys[60].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__stu__valid        ( PeArray2Sys[61].pe__stu__valid             ),      
        .pe61__stu__cntl         ( PeArray2Sys[61].pe__stu__cntl              ),      
        .stu__pe61__ready        ( 1'b1     ),      
        //.stu__pe61__ready        ( PeArray2Sys[61].cb_test.stu__pe__ready     ),      
        .pe61__stu__type         ( PeArray2Sys[61].pe__stu__type              ),      
        .pe61__stu__data         ( PeArray2Sys[61].pe__stu__data              ),      
        .pe61__stu__oob_data     ( PeArray2Sys[61].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__stu__valid        ( PeArray2Sys[62].pe__stu__valid             ),      
        .pe62__stu__cntl         ( PeArray2Sys[62].pe__stu__cntl              ),      
        .stu__pe62__ready        ( 1'b1     ),      
        //.stu__pe62__ready        ( PeArray2Sys[62].cb_test.stu__pe__ready     ),      
        .pe62__stu__type         ( PeArray2Sys[62].pe__stu__type              ),      
        .pe62__stu__data         ( PeArray2Sys[62].pe__stu__data              ),      
        .pe62__stu__oob_data     ( PeArray2Sys[62].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__stu__valid        ( PeArray2Sys[63].pe__stu__valid             ),      
        .pe63__stu__cntl         ( PeArray2Sys[63].pe__stu__cntl              ),      
        .stu__pe63__ready        ( 1'b1     ),      
        //.stu__pe63__ready        ( PeArray2Sys[63].cb_test.stu__pe__ready     ),      
        .pe63__stu__type         ( PeArray2Sys[63].pe__stu__type              ),      
        .pe63__stu__data         ( PeArray2Sys[63].pe__stu__data              ),      
        .pe63__stu__oob_data     ( PeArray2Sys[63].pe__stu__oob_data          ),      
        