
    input                                          pe0__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe0__stu__cntl           ;
    output                                         stu__pe0__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe0__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe0__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe0__stu__oob_data       ;

    input                                          pe1__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe1__stu__cntl           ;
    output                                         stu__pe1__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe1__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe1__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe1__stu__oob_data       ;

    input                                          pe2__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe2__stu__cntl           ;
    output                                         stu__pe2__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe2__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe2__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe2__stu__oob_data       ;

    input                                          pe3__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe3__stu__cntl           ;
    output                                         stu__pe3__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe3__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe3__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe3__stu__oob_data       ;

    input                                          pe4__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe4__stu__cntl           ;
    output                                         stu__pe4__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe4__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe4__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe4__stu__oob_data       ;

    input                                          pe5__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe5__stu__cntl           ;
    output                                         stu__pe5__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe5__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe5__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe5__stu__oob_data       ;

    input                                          pe6__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe6__stu__cntl           ;
    output                                         stu__pe6__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe6__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe6__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe6__stu__oob_data       ;

    input                                          pe7__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe7__stu__cntl           ;
    output                                         stu__pe7__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe7__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe7__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe7__stu__oob_data       ;

    input                                          pe8__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe8__stu__cntl           ;
    output                                         stu__pe8__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe8__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe8__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe8__stu__oob_data       ;

    input                                          pe9__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe9__stu__cntl           ;
    output                                         stu__pe9__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe9__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe9__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe9__stu__oob_data       ;

    input                                          pe10__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe10__stu__cntl           ;
    output                                         stu__pe10__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe10__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe10__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe10__stu__oob_data       ;

    input                                          pe11__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe11__stu__cntl           ;
    output                                         stu__pe11__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe11__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe11__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe11__stu__oob_data       ;

    input                                          pe12__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe12__stu__cntl           ;
    output                                         stu__pe12__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe12__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe12__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe12__stu__oob_data       ;

    input                                          pe13__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe13__stu__cntl           ;
    output                                         stu__pe13__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe13__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe13__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe13__stu__oob_data       ;

    input                                          pe14__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe14__stu__cntl           ;
    output                                         stu__pe14__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe14__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe14__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe14__stu__oob_data       ;

    input                                          pe15__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe15__stu__cntl           ;
    output                                         stu__pe15__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe15__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe15__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe15__stu__oob_data       ;

    input                                          pe16__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe16__stu__cntl           ;
    output                                         stu__pe16__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe16__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe16__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe16__stu__oob_data       ;

    input                                          pe17__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe17__stu__cntl           ;
    output                                         stu__pe17__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe17__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe17__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe17__stu__oob_data       ;

    input                                          pe18__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe18__stu__cntl           ;
    output                                         stu__pe18__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe18__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe18__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe18__stu__oob_data       ;

    input                                          pe19__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe19__stu__cntl           ;
    output                                         stu__pe19__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe19__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe19__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe19__stu__oob_data       ;

    input                                          pe20__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe20__stu__cntl           ;
    output                                         stu__pe20__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe20__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe20__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe20__stu__oob_data       ;

    input                                          pe21__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe21__stu__cntl           ;
    output                                         stu__pe21__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe21__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe21__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe21__stu__oob_data       ;

    input                                          pe22__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe22__stu__cntl           ;
    output                                         stu__pe22__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe22__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe22__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe22__stu__oob_data       ;

    input                                          pe23__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe23__stu__cntl           ;
    output                                         stu__pe23__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe23__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe23__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe23__stu__oob_data       ;

    input                                          pe24__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe24__stu__cntl           ;
    output                                         stu__pe24__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe24__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe24__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe24__stu__oob_data       ;

    input                                          pe25__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe25__stu__cntl           ;
    output                                         stu__pe25__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe25__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe25__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe25__stu__oob_data       ;

    input                                          pe26__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe26__stu__cntl           ;
    output                                         stu__pe26__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe26__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe26__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe26__stu__oob_data       ;

    input                                          pe27__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe27__stu__cntl           ;
    output                                         stu__pe27__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe27__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe27__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe27__stu__oob_data       ;

    input                                          pe28__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe28__stu__cntl           ;
    output                                         stu__pe28__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe28__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe28__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe28__stu__oob_data       ;

    input                                          pe29__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe29__stu__cntl           ;
    output                                         stu__pe29__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe29__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe29__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe29__stu__oob_data       ;

    input                                          pe30__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe30__stu__cntl           ;
    output                                         stu__pe30__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe30__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe30__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe30__stu__oob_data       ;

    input                                          pe31__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe31__stu__cntl           ;
    output                                         stu__pe31__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe31__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe31__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe31__stu__oob_data       ;

    input                                          pe32__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe32__stu__cntl           ;
    output                                         stu__pe32__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe32__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe32__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe32__stu__oob_data       ;

    input                                          pe33__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe33__stu__cntl           ;
    output                                         stu__pe33__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe33__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe33__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe33__stu__oob_data       ;

    input                                          pe34__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe34__stu__cntl           ;
    output                                         stu__pe34__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe34__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe34__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe34__stu__oob_data       ;

    input                                          pe35__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe35__stu__cntl           ;
    output                                         stu__pe35__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe35__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe35__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe35__stu__oob_data       ;

    input                                          pe36__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe36__stu__cntl           ;
    output                                         stu__pe36__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe36__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe36__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe36__stu__oob_data       ;

    input                                          pe37__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe37__stu__cntl           ;
    output                                         stu__pe37__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe37__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe37__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe37__stu__oob_data       ;

    input                                          pe38__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe38__stu__cntl           ;
    output                                         stu__pe38__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe38__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe38__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe38__stu__oob_data       ;

    input                                          pe39__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe39__stu__cntl           ;
    output                                         stu__pe39__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe39__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe39__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe39__stu__oob_data       ;

    input                                          pe40__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe40__stu__cntl           ;
    output                                         stu__pe40__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe40__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe40__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe40__stu__oob_data       ;

    input                                          pe41__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe41__stu__cntl           ;
    output                                         stu__pe41__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe41__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe41__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe41__stu__oob_data       ;

    input                                          pe42__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe42__stu__cntl           ;
    output                                         stu__pe42__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe42__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe42__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe42__stu__oob_data       ;

    input                                          pe43__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe43__stu__cntl           ;
    output                                         stu__pe43__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe43__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe43__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe43__stu__oob_data       ;

    input                                          pe44__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe44__stu__cntl           ;
    output                                         stu__pe44__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe44__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe44__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe44__stu__oob_data       ;

    input                                          pe45__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe45__stu__cntl           ;
    output                                         stu__pe45__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe45__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe45__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe45__stu__oob_data       ;

    input                                          pe46__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe46__stu__cntl           ;
    output                                         stu__pe46__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe46__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe46__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe46__stu__oob_data       ;

    input                                          pe47__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe47__stu__cntl           ;
    output                                         stu__pe47__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe47__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe47__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe47__stu__oob_data       ;

    input                                          pe48__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe48__stu__cntl           ;
    output                                         stu__pe48__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe48__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe48__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe48__stu__oob_data       ;

    input                                          pe49__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe49__stu__cntl           ;
    output                                         stu__pe49__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe49__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe49__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe49__stu__oob_data       ;

    input                                          pe50__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe50__stu__cntl           ;
    output                                         stu__pe50__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe50__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe50__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe50__stu__oob_data       ;

    input                                          pe51__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe51__stu__cntl           ;
    output                                         stu__pe51__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe51__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe51__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe51__stu__oob_data       ;

    input                                          pe52__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe52__stu__cntl           ;
    output                                         stu__pe52__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe52__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe52__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe52__stu__oob_data       ;

    input                                          pe53__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe53__stu__cntl           ;
    output                                         stu__pe53__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe53__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe53__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe53__stu__oob_data       ;

    input                                          pe54__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe54__stu__cntl           ;
    output                                         stu__pe54__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe54__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe54__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe54__stu__oob_data       ;

    input                                          pe55__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe55__stu__cntl           ;
    output                                         stu__pe55__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe55__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe55__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe55__stu__oob_data       ;

    input                                          pe56__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe56__stu__cntl           ;
    output                                         stu__pe56__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe56__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe56__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe56__stu__oob_data       ;

    input                                          pe57__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe57__stu__cntl           ;
    output                                         stu__pe57__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe57__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe57__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe57__stu__oob_data       ;

    input                                          pe58__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe58__stu__cntl           ;
    output                                         stu__pe58__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe58__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe58__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe58__stu__oob_data       ;

    input                                          pe59__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe59__stu__cntl           ;
    output                                         stu__pe59__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe59__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe59__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe59__stu__oob_data       ;

    input                                          pe60__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe60__stu__cntl           ;
    output                                         stu__pe60__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe60__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe60__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe60__stu__oob_data       ;

    input                                          pe61__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe61__stu__cntl           ;
    output                                         stu__pe61__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe61__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe61__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe61__stu__oob_data       ;

    input                                          pe62__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe62__stu__cntl           ;
    output                                         stu__pe62__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe62__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe62__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe62__stu__oob_data       ;

    input                                          pe63__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe63__stu__cntl           ;
    output                                         stu__pe63__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe63__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe63__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe63__stu__oob_data       ;

