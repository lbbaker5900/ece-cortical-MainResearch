
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr0__std__oob_cntl            ;
  output                                          mgr0__std__oob_valid           ;
  input                                           std__mgr0__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr0__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr0__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr1__std__oob_cntl            ;
  output                                          mgr1__std__oob_valid           ;
  input                                           std__mgr1__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr1__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr1__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr2__std__oob_cntl            ;
  output                                          mgr2__std__oob_valid           ;
  input                                           std__mgr2__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr2__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr2__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr3__std__oob_cntl            ;
  output                                          mgr3__std__oob_valid           ;
  input                                           std__mgr3__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr3__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr3__std__oob_data            ;