
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[0].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[0].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[0].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[0].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[0].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[0].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[1].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[1].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[1].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[1].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[1].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[1].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[2].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[2].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[2].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[2].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[2].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[2].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[3].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[3].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[3].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[3].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[3].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[3].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[4].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[4].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[4].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[4].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[4].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[4].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[4].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[5].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[5].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[5].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[5].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[5].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[5].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[5].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[6].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[6].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[6].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[6].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[6].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[6].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[6].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[7].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[7].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[7].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[7].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[7].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[7].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[7].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[8].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[8].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[8].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[8].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[8].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[8].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[8].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[9].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[9].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[9].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[9].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[9].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[9].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[9].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[10].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[10].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[10].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[10].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[10].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[10].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[10].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[11].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[11].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[11].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[11].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[11].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[11].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[11].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[12].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[12].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[12].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[12].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[12].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[12].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[12].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[13].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[13].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[13].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[13].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[13].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[13].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[13].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[14].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[14].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[14].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[14].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[14].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[14].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[14].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[15].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[15].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[15].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[15].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[15].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[15].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[15].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[16].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[16].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[16].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[16].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[16].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[16].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[16].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[17].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[17].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[17].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[17].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[17].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[17].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[17].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[18].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[18].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[18].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[18].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[18].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[18].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[18].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[19].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[19].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[19].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[19].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[19].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[19].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[19].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[20].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[20].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[20].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[20].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[20].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[20].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[20].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[21].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[21].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[21].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[21].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[21].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[21].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[21].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[22].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[22].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[22].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[22].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[22].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[22].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[22].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[23].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[23].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[23].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[23].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[23].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[23].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[23].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[24].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[24].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[24].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[24].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[24].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[24].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[24].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[25].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[25].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[25].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[25].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[25].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[25].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[25].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[26].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[26].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[26].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[26].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[26].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[26].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[26].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[27].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[27].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[27].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[27].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[27].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[27].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[27].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[28].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[28].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[28].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[28].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[28].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[28].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[28].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[29].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[29].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[29].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[29].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[29].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[29].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[29].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[30].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[30].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[30].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[30].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[30].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[30].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[30].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[31].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[31].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[31].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[31].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[31].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[31].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[31].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[32].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[32].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[32].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[32].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[32].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[32].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[32].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[33].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[33].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[33].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[33].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[33].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[33].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[33].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[34].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[34].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[34].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[34].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[34].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[34].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[34].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[35].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[35].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[35].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[35].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[35].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[35].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[35].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[36].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[36].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[36].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[36].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[36].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[36].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[36].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[37].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[37].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[37].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[37].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[37].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[37].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[37].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[38].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[38].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[38].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[38].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[38].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[38].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[38].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[39].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[39].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[39].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[39].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[39].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[39].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[39].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[40].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[40].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[40].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[40].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[40].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[40].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[40].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[41].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[41].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[41].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[41].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[41].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[41].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[41].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[42].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[42].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[42].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[42].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[42].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[42].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[42].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[43].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[43].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[43].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[43].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[43].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[43].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[43].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[44].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[44].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[44].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[44].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[44].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[44].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[44].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[45].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[45].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[45].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[45].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[45].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[45].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[45].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[46].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[46].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[46].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[46].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[46].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[46].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[46].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[47].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[47].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[47].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[47].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[47].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[47].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[47].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[48].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[48].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[48].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[48].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[48].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[48].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[48].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[49].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[49].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[49].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[49].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[49].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[49].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[49].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[50].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[50].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[50].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[50].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[50].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[50].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[50].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[51].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[51].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[51].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[51].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[51].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[51].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[51].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[52].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[52].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[52].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[52].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[52].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[52].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[52].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[53].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[53].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[53].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[53].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[53].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[53].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[53].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[54].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[54].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[54].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[54].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[54].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[54].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[54].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[55].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[55].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[55].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[55].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[55].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[55].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[55].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[56].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[56].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[56].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[56].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[56].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[56].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[56].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[57].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[57].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[57].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[57].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[57].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[57].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[57].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[58].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[58].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[58].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[58].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[58].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[58].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[58].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[59].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[59].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[59].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[59].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[59].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[59].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[59].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[60].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[60].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[60].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[60].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[60].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[60].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[60].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[61].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[61].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[61].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[61].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[61].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[61].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[61].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[62].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[62].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[62].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[62].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[62].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[62].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[62].pe.ldst__memc__read_valid  = 1'b0; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane0_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane0_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane0_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane0_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane0_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane0_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane0_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane0_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane1_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane1_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane1_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane1_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane1_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane1_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane1_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane1_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane2_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane2_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane2_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane2_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane2_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane2_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane2_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane2_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane3_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane3_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane3_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane3_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane3_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane3_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane3_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane3_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane4_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane4_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane4_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane4_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane4_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane4_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane4_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane4_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane5_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane5_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane5_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane5_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane5_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane5_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane5_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane5_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane6_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane6_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane6_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane6_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane6_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane6_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane6_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane6_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane7_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane7_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane7_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane7_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane7_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane7_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane7_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane7_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane8_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane8_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane8_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane8_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane8_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane8_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane8_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane8_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane9_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane9_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane9_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane9_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane9_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane9_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane9_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane9_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane10_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane10_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane10_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane10_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane10_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane10_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane10_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane10_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane11_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane11_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane11_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane11_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane11_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane11_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane11_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane11_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane12_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane12_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane12_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane12_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane12_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane12_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane12_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane12_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane13_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane13_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane13_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane13_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane13_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane13_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane13_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane13_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane14_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane14_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane14_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane14_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane14_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane14_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane14_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane14_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane15_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane15_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane15_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane15_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane15_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane15_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane15_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane15_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane16_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane16_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane16_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane16_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane16_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane16_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane16_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane16_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane17_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane17_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane17_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane17_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane17_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane17_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane17_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane17_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane18_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane18_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane18_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane18_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane18_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane18_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane18_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane18_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane19_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane19_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane19_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane19_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane19_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane19_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane19_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane19_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane20_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane20_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane20_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane20_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane20_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane20_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane20_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane20_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane21_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane21_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane21_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane21_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane21_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane21_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane21_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane21_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane22_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane22_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane22_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane22_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane22_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane22_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane22_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane22_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane23_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane23_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane23_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane23_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane23_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane23_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane23_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane23_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane24_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane24_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane24_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane24_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane24_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane24_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane24_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane24_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane25_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane25_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane25_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane25_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane25_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane25_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane25_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane25_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane26_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane26_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane26_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane26_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane26_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane26_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane26_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane26_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane27_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane27_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane27_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane27_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane27_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane27_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane27_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane27_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane28_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane28_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane28_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane28_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane28_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane28_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane28_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane28_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane29_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane29_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane29_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane29_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane29_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane29_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane29_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane29_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane30_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane30_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane30_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane30_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane30_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane30_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane30_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane30_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane31_r128 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane31_r129 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane31_r130 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane31_r131 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane31_r132 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane31_r133 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane31_r134 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane31_r135 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[63].pe.ldst__memc__request   = 1'b0 ; 
    force pe_array_inst.pe_inst[63].pe.ldst__memc__released  = 1'b1 ; 
    force pe_array_inst.pe_inst[63].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[63].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[63].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[63].pe.ldst__memc__write_valid = 1'b0; 
    force pe_array_inst.pe_inst[63].pe.ldst__memc__read_valid  = 1'b0; 