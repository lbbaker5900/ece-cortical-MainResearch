
  wire  sys__pe__allSynchronized = pe_inst[0].pe__sys__thisSynchronized & 
                                   pe_inst[1].pe__sys__thisSynchronized & 
                                   pe_inst[2].pe__sys__thisSynchronized & 
                                   pe_inst[3].pe__sys__thisSynchronized & 
                                   pe_inst[4].pe__sys__thisSynchronized & 
                                   pe_inst[5].pe__sys__thisSynchronized & 
                                   pe_inst[6].pe__sys__thisSynchronized & 
                                   pe_inst[7].pe__sys__thisSynchronized & 
                                   pe_inst[8].pe__sys__thisSynchronized & 
                                   pe_inst[9].pe__sys__thisSynchronized & 
                                   pe_inst[10].pe__sys__thisSynchronized & 
                                   pe_inst[11].pe__sys__thisSynchronized & 
                                   pe_inst[12].pe__sys__thisSynchronized & 
                                   pe_inst[13].pe__sys__thisSynchronized & 
                                   pe_inst[14].pe__sys__thisSynchronized & 
                                   pe_inst[15].pe__sys__thisSynchronized & 
                                   pe_inst[16].pe__sys__thisSynchronized & 
                                   pe_inst[17].pe__sys__thisSynchronized & 
                                   pe_inst[18].pe__sys__thisSynchronized & 
                                   pe_inst[19].pe__sys__thisSynchronized & 
                                   pe_inst[20].pe__sys__thisSynchronized & 
                                   pe_inst[21].pe__sys__thisSynchronized & 
                                   pe_inst[22].pe__sys__thisSynchronized & 
                                   pe_inst[23].pe__sys__thisSynchronized & 
                                   pe_inst[24].pe__sys__thisSynchronized & 
                                   pe_inst[25].pe__sys__thisSynchronized & 
                                   pe_inst[26].pe__sys__thisSynchronized & 
                                   pe_inst[27].pe__sys__thisSynchronized & 
                                   pe_inst[28].pe__sys__thisSynchronized & 
                                   pe_inst[29].pe__sys__thisSynchronized & 
                                   pe_inst[30].pe__sys__thisSynchronized & 
                                   pe_inst[31].pe__sys__thisSynchronized & 
                                   pe_inst[32].pe__sys__thisSynchronized & 
                                   pe_inst[33].pe__sys__thisSynchronized & 
                                   pe_inst[34].pe__sys__thisSynchronized & 
                                   pe_inst[35].pe__sys__thisSynchronized & 
                                   pe_inst[36].pe__sys__thisSynchronized & 
                                   pe_inst[37].pe__sys__thisSynchronized & 
                                   pe_inst[38].pe__sys__thisSynchronized & 
                                   pe_inst[39].pe__sys__thisSynchronized & 
                                   pe_inst[40].pe__sys__thisSynchronized & 
                                   pe_inst[41].pe__sys__thisSynchronized & 
                                   pe_inst[42].pe__sys__thisSynchronized & 
                                   pe_inst[43].pe__sys__thisSynchronized & 
                                   pe_inst[44].pe__sys__thisSynchronized & 
                                   pe_inst[45].pe__sys__thisSynchronized & 
                                   pe_inst[46].pe__sys__thisSynchronized & 
                                   pe_inst[47].pe__sys__thisSynchronized & 
                                   pe_inst[48].pe__sys__thisSynchronized & 
                                   pe_inst[49].pe__sys__thisSynchronized & 
                                   pe_inst[50].pe__sys__thisSynchronized & 
                                   pe_inst[51].pe__sys__thisSynchronized & 
                                   pe_inst[52].pe__sys__thisSynchronized & 
                                   pe_inst[53].pe__sys__thisSynchronized & 
                                   pe_inst[54].pe__sys__thisSynchronized & 
                                   pe_inst[55].pe__sys__thisSynchronized & 
                                   pe_inst[56].pe__sys__thisSynchronized & 
                                   pe_inst[57].pe__sys__thisSynchronized & 
                                   pe_inst[58].pe__sys__thisSynchronized & 
                                   pe_inst[59].pe__sys__thisSynchronized & 
                                   pe_inst[60].pe__sys__thisSynchronized & 
                                   pe_inst[61].pe__sys__thisSynchronized & 
                                   pe_inst[62].pe__sys__thisSynchronized & 
                                   pe_inst[63].pe__sys__thisSynchronized ; 