
        // PE 0, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane0_strm0_ready         ( DownstreamStackBusLane[0][0].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane0_strm0_cntl          ( DownstreamStackBusLane[0][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane0_strm0_data          ( DownstreamStackBusLane[0][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane0_strm0_data_valid    ( DownstreamStackBusLane[0][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane0_strm1_ready         ( DownstreamStackBusLane[0][0].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane0_strm1_cntl          ( DownstreamStackBusLane[0][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane0_strm1_data          ( DownstreamStackBusLane[0][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane0_strm1_data_valid    ( DownstreamStackBusLane[0][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane1_strm0_ready         ( DownstreamStackBusLane[0][1].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane1_strm0_cntl          ( DownstreamStackBusLane[0][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane1_strm0_data          ( DownstreamStackBusLane[0][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane1_strm0_data_valid    ( DownstreamStackBusLane[0][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane1_strm1_ready         ( DownstreamStackBusLane[0][1].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane1_strm1_cntl          ( DownstreamStackBusLane[0][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane1_strm1_data          ( DownstreamStackBusLane[0][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane1_strm1_data_valid    ( DownstreamStackBusLane[0][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane2_strm0_ready         ( DownstreamStackBusLane[0][2].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane2_strm0_cntl          ( DownstreamStackBusLane[0][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane2_strm0_data          ( DownstreamStackBusLane[0][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane2_strm0_data_valid    ( DownstreamStackBusLane[0][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane2_strm1_ready         ( DownstreamStackBusLane[0][2].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane2_strm1_cntl          ( DownstreamStackBusLane[0][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane2_strm1_data          ( DownstreamStackBusLane[0][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane2_strm1_data_valid    ( DownstreamStackBusLane[0][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane3_strm0_ready         ( DownstreamStackBusLane[0][3].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane3_strm0_cntl          ( DownstreamStackBusLane[0][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane3_strm0_data          ( DownstreamStackBusLane[0][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane3_strm0_data_valid    ( DownstreamStackBusLane[0][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane3_strm1_ready         ( DownstreamStackBusLane[0][3].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane3_strm1_cntl          ( DownstreamStackBusLane[0][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane3_strm1_data          ( DownstreamStackBusLane[0][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane3_strm1_data_valid    ( DownstreamStackBusLane[0][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane4_strm0_ready         ( DownstreamStackBusLane[0][4].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane4_strm0_cntl          ( DownstreamStackBusLane[0][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane4_strm0_data          ( DownstreamStackBusLane[0][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane4_strm0_data_valid    ( DownstreamStackBusLane[0][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane4_strm1_ready         ( DownstreamStackBusLane[0][4].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane4_strm1_cntl          ( DownstreamStackBusLane[0][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane4_strm1_data          ( DownstreamStackBusLane[0][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane4_strm1_data_valid    ( DownstreamStackBusLane[0][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane5_strm0_ready         ( DownstreamStackBusLane[0][5].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane5_strm0_cntl          ( DownstreamStackBusLane[0][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane5_strm0_data          ( DownstreamStackBusLane[0][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane5_strm0_data_valid    ( DownstreamStackBusLane[0][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane5_strm1_ready         ( DownstreamStackBusLane[0][5].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane5_strm1_cntl          ( DownstreamStackBusLane[0][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane5_strm1_data          ( DownstreamStackBusLane[0][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane5_strm1_data_valid    ( DownstreamStackBusLane[0][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane6_strm0_ready         ( DownstreamStackBusLane[0][6].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane6_strm0_cntl          ( DownstreamStackBusLane[0][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane6_strm0_data          ( DownstreamStackBusLane[0][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane6_strm0_data_valid    ( DownstreamStackBusLane[0][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane6_strm1_ready         ( DownstreamStackBusLane[0][6].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane6_strm1_cntl          ( DownstreamStackBusLane[0][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane6_strm1_data          ( DownstreamStackBusLane[0][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane6_strm1_data_valid    ( DownstreamStackBusLane[0][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane7_strm0_ready         ( DownstreamStackBusLane[0][7].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane7_strm0_cntl          ( DownstreamStackBusLane[0][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane7_strm0_data          ( DownstreamStackBusLane[0][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane7_strm0_data_valid    ( DownstreamStackBusLane[0][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane7_strm1_ready         ( DownstreamStackBusLane[0][7].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane7_strm1_cntl          ( DownstreamStackBusLane[0][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane7_strm1_data          ( DownstreamStackBusLane[0][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane7_strm1_data_valid    ( DownstreamStackBusLane[0][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane8_strm0_ready         ( DownstreamStackBusLane[0][8].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane8_strm0_cntl          ( DownstreamStackBusLane[0][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane8_strm0_data          ( DownstreamStackBusLane[0][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane8_strm0_data_valid    ( DownstreamStackBusLane[0][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane8_strm1_ready         ( DownstreamStackBusLane[0][8].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane8_strm1_cntl          ( DownstreamStackBusLane[0][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane8_strm1_data          ( DownstreamStackBusLane[0][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane8_strm1_data_valid    ( DownstreamStackBusLane[0][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane9_strm0_ready         ( DownstreamStackBusLane[0][9].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane9_strm0_cntl          ( DownstreamStackBusLane[0][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane9_strm0_data          ( DownstreamStackBusLane[0][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane9_strm0_data_valid    ( DownstreamStackBusLane[0][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane9_strm1_ready         ( DownstreamStackBusLane[0][9].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane9_strm1_cntl          ( DownstreamStackBusLane[0][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane9_strm1_data          ( DownstreamStackBusLane[0][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane9_strm1_data_valid    ( DownstreamStackBusLane[0][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane10_strm0_ready         ( DownstreamStackBusLane[0][10].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane10_strm0_cntl          ( DownstreamStackBusLane[0][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane10_strm0_data          ( DownstreamStackBusLane[0][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane10_strm0_data_valid    ( DownstreamStackBusLane[0][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane10_strm1_ready         ( DownstreamStackBusLane[0][10].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane10_strm1_cntl          ( DownstreamStackBusLane[0][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane10_strm1_data          ( DownstreamStackBusLane[0][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane10_strm1_data_valid    ( DownstreamStackBusLane[0][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane11_strm0_ready         ( DownstreamStackBusLane[0][11].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane11_strm0_cntl          ( DownstreamStackBusLane[0][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane11_strm0_data          ( DownstreamStackBusLane[0][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane11_strm0_data_valid    ( DownstreamStackBusLane[0][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane11_strm1_ready         ( DownstreamStackBusLane[0][11].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane11_strm1_cntl          ( DownstreamStackBusLane[0][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane11_strm1_data          ( DownstreamStackBusLane[0][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane11_strm1_data_valid    ( DownstreamStackBusLane[0][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane12_strm0_ready         ( DownstreamStackBusLane[0][12].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane12_strm0_cntl          ( DownstreamStackBusLane[0][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane12_strm0_data          ( DownstreamStackBusLane[0][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane12_strm0_data_valid    ( DownstreamStackBusLane[0][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane12_strm1_ready         ( DownstreamStackBusLane[0][12].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane12_strm1_cntl          ( DownstreamStackBusLane[0][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane12_strm1_data          ( DownstreamStackBusLane[0][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane12_strm1_data_valid    ( DownstreamStackBusLane[0][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane13_strm0_ready         ( DownstreamStackBusLane[0][13].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane13_strm0_cntl          ( DownstreamStackBusLane[0][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane13_strm0_data          ( DownstreamStackBusLane[0][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane13_strm0_data_valid    ( DownstreamStackBusLane[0][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane13_strm1_ready         ( DownstreamStackBusLane[0][13].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane13_strm1_cntl          ( DownstreamStackBusLane[0][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane13_strm1_data          ( DownstreamStackBusLane[0][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane13_strm1_data_valid    ( DownstreamStackBusLane[0][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane14_strm0_ready         ( DownstreamStackBusLane[0][14].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane14_strm0_cntl          ( DownstreamStackBusLane[0][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane14_strm0_data          ( DownstreamStackBusLane[0][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane14_strm0_data_valid    ( DownstreamStackBusLane[0][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane14_strm1_ready         ( DownstreamStackBusLane[0][14].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane14_strm1_cntl          ( DownstreamStackBusLane[0][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane14_strm1_data          ( DownstreamStackBusLane[0][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane14_strm1_data_valid    ( DownstreamStackBusLane[0][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane15_strm0_ready         ( DownstreamStackBusLane[0][15].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane15_strm0_cntl          ( DownstreamStackBusLane[0][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane15_strm0_data          ( DownstreamStackBusLane[0][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane15_strm0_data_valid    ( DownstreamStackBusLane[0][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane15_strm1_ready         ( DownstreamStackBusLane[0][15].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane15_strm1_cntl          ( DownstreamStackBusLane[0][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane15_strm1_data          ( DownstreamStackBusLane[0][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane15_strm1_data_valid    ( DownstreamStackBusLane[0][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane16_strm0_ready         ( DownstreamStackBusLane[0][16].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane16_strm0_cntl          ( DownstreamStackBusLane[0][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane16_strm0_data          ( DownstreamStackBusLane[0][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane16_strm0_data_valid    ( DownstreamStackBusLane[0][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane16_strm1_ready         ( DownstreamStackBusLane[0][16].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane16_strm1_cntl          ( DownstreamStackBusLane[0][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane16_strm1_data          ( DownstreamStackBusLane[0][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane16_strm1_data_valid    ( DownstreamStackBusLane[0][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane17_strm0_ready         ( DownstreamStackBusLane[0][17].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane17_strm0_cntl          ( DownstreamStackBusLane[0][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane17_strm0_data          ( DownstreamStackBusLane[0][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane17_strm0_data_valid    ( DownstreamStackBusLane[0][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane17_strm1_ready         ( DownstreamStackBusLane[0][17].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane17_strm1_cntl          ( DownstreamStackBusLane[0][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane17_strm1_data          ( DownstreamStackBusLane[0][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane17_strm1_data_valid    ( DownstreamStackBusLane[0][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane18_strm0_ready         ( DownstreamStackBusLane[0][18].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane18_strm0_cntl          ( DownstreamStackBusLane[0][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane18_strm0_data          ( DownstreamStackBusLane[0][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane18_strm0_data_valid    ( DownstreamStackBusLane[0][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane18_strm1_ready         ( DownstreamStackBusLane[0][18].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane18_strm1_cntl          ( DownstreamStackBusLane[0][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane18_strm1_data          ( DownstreamStackBusLane[0][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane18_strm1_data_valid    ( DownstreamStackBusLane[0][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane19_strm0_ready         ( DownstreamStackBusLane[0][19].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane19_strm0_cntl          ( DownstreamStackBusLane[0][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane19_strm0_data          ( DownstreamStackBusLane[0][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane19_strm0_data_valid    ( DownstreamStackBusLane[0][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane19_strm1_ready         ( DownstreamStackBusLane[0][19].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane19_strm1_cntl          ( DownstreamStackBusLane[0][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane19_strm1_data          ( DownstreamStackBusLane[0][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane19_strm1_data_valid    ( DownstreamStackBusLane[0][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane20_strm0_ready         ( DownstreamStackBusLane[0][20].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane20_strm0_cntl          ( DownstreamStackBusLane[0][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane20_strm0_data          ( DownstreamStackBusLane[0][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane20_strm0_data_valid    ( DownstreamStackBusLane[0][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane20_strm1_ready         ( DownstreamStackBusLane[0][20].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane20_strm1_cntl          ( DownstreamStackBusLane[0][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane20_strm1_data          ( DownstreamStackBusLane[0][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane20_strm1_data_valid    ( DownstreamStackBusLane[0][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane21_strm0_ready         ( DownstreamStackBusLane[0][21].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane21_strm0_cntl          ( DownstreamStackBusLane[0][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane21_strm0_data          ( DownstreamStackBusLane[0][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane21_strm0_data_valid    ( DownstreamStackBusLane[0][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane21_strm1_ready         ( DownstreamStackBusLane[0][21].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane21_strm1_cntl          ( DownstreamStackBusLane[0][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane21_strm1_data          ( DownstreamStackBusLane[0][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane21_strm1_data_valid    ( DownstreamStackBusLane[0][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane22_strm0_ready         ( DownstreamStackBusLane[0][22].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane22_strm0_cntl          ( DownstreamStackBusLane[0][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane22_strm0_data          ( DownstreamStackBusLane[0][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane22_strm0_data_valid    ( DownstreamStackBusLane[0][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane22_strm1_ready         ( DownstreamStackBusLane[0][22].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane22_strm1_cntl          ( DownstreamStackBusLane[0][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane22_strm1_data          ( DownstreamStackBusLane[0][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane22_strm1_data_valid    ( DownstreamStackBusLane[0][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane23_strm0_ready         ( DownstreamStackBusLane[0][23].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane23_strm0_cntl          ( DownstreamStackBusLane[0][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane23_strm0_data          ( DownstreamStackBusLane[0][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane23_strm0_data_valid    ( DownstreamStackBusLane[0][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane23_strm1_ready         ( DownstreamStackBusLane[0][23].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane23_strm1_cntl          ( DownstreamStackBusLane[0][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane23_strm1_data          ( DownstreamStackBusLane[0][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane23_strm1_data_valid    ( DownstreamStackBusLane[0][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane24_strm0_ready         ( DownstreamStackBusLane[0][24].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane24_strm0_cntl          ( DownstreamStackBusLane[0][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane24_strm0_data          ( DownstreamStackBusLane[0][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane24_strm0_data_valid    ( DownstreamStackBusLane[0][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane24_strm1_ready         ( DownstreamStackBusLane[0][24].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane24_strm1_cntl          ( DownstreamStackBusLane[0][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane24_strm1_data          ( DownstreamStackBusLane[0][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane24_strm1_data_valid    ( DownstreamStackBusLane[0][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane25_strm0_ready         ( DownstreamStackBusLane[0][25].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane25_strm0_cntl          ( DownstreamStackBusLane[0][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane25_strm0_data          ( DownstreamStackBusLane[0][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane25_strm0_data_valid    ( DownstreamStackBusLane[0][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane25_strm1_ready         ( DownstreamStackBusLane[0][25].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane25_strm1_cntl          ( DownstreamStackBusLane[0][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane25_strm1_data          ( DownstreamStackBusLane[0][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane25_strm1_data_valid    ( DownstreamStackBusLane[0][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane26_strm0_ready         ( DownstreamStackBusLane[0][26].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane26_strm0_cntl          ( DownstreamStackBusLane[0][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane26_strm0_data          ( DownstreamStackBusLane[0][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane26_strm0_data_valid    ( DownstreamStackBusLane[0][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane26_strm1_ready         ( DownstreamStackBusLane[0][26].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane26_strm1_cntl          ( DownstreamStackBusLane[0][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane26_strm1_data          ( DownstreamStackBusLane[0][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane26_strm1_data_valid    ( DownstreamStackBusLane[0][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane27_strm0_ready         ( DownstreamStackBusLane[0][27].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane27_strm0_cntl          ( DownstreamStackBusLane[0][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane27_strm0_data          ( DownstreamStackBusLane[0][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane27_strm0_data_valid    ( DownstreamStackBusLane[0][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane27_strm1_ready         ( DownstreamStackBusLane[0][27].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane27_strm1_cntl          ( DownstreamStackBusLane[0][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane27_strm1_data          ( DownstreamStackBusLane[0][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane27_strm1_data_valid    ( DownstreamStackBusLane[0][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane28_strm0_ready         ( DownstreamStackBusLane[0][28].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane28_strm0_cntl          ( DownstreamStackBusLane[0][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane28_strm0_data          ( DownstreamStackBusLane[0][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane28_strm0_data_valid    ( DownstreamStackBusLane[0][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane28_strm1_ready         ( DownstreamStackBusLane[0][28].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane28_strm1_cntl          ( DownstreamStackBusLane[0][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane28_strm1_data          ( DownstreamStackBusLane[0][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane28_strm1_data_valid    ( DownstreamStackBusLane[0][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane29_strm0_ready         ( DownstreamStackBusLane[0][29].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane29_strm0_cntl          ( DownstreamStackBusLane[0][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane29_strm0_data          ( DownstreamStackBusLane[0][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane29_strm0_data_valid    ( DownstreamStackBusLane[0][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane29_strm1_ready         ( DownstreamStackBusLane[0][29].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane29_strm1_cntl          ( DownstreamStackBusLane[0][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane29_strm1_data          ( DownstreamStackBusLane[0][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane29_strm1_data_valid    ( DownstreamStackBusLane[0][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane30_strm0_ready         ( DownstreamStackBusLane[0][30].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane30_strm0_cntl          ( DownstreamStackBusLane[0][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane30_strm0_data          ( DownstreamStackBusLane[0][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane30_strm0_data_valid    ( DownstreamStackBusLane[0][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane30_strm1_ready         ( DownstreamStackBusLane[0][30].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane30_strm1_cntl          ( DownstreamStackBusLane[0][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane30_strm1_data          ( DownstreamStackBusLane[0][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane30_strm1_data_valid    ( DownstreamStackBusLane[0][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane31_strm0_ready         ( DownstreamStackBusLane[0][31].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane31_strm0_cntl          ( DownstreamStackBusLane[0][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane31_strm0_data          ( DownstreamStackBusLane[0][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane31_strm0_data_valid    ( DownstreamStackBusLane[0][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane31_strm1_ready         ( DownstreamStackBusLane[0][31].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane31_strm1_cntl          ( DownstreamStackBusLane[0][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane31_strm1_data          ( DownstreamStackBusLane[0][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane31_strm1_data_valid    ( DownstreamStackBusLane[0][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane0_strm0_ready         ( DownstreamStackBusLane[1][0].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane0_strm0_cntl          ( DownstreamStackBusLane[1][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane0_strm0_data          ( DownstreamStackBusLane[1][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane0_strm0_data_valid    ( DownstreamStackBusLane[1][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane0_strm1_ready         ( DownstreamStackBusLane[1][0].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane0_strm1_cntl          ( DownstreamStackBusLane[1][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane0_strm1_data          ( DownstreamStackBusLane[1][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane0_strm1_data_valid    ( DownstreamStackBusLane[1][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane1_strm0_ready         ( DownstreamStackBusLane[1][1].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane1_strm0_cntl          ( DownstreamStackBusLane[1][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane1_strm0_data          ( DownstreamStackBusLane[1][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane1_strm0_data_valid    ( DownstreamStackBusLane[1][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane1_strm1_ready         ( DownstreamStackBusLane[1][1].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane1_strm1_cntl          ( DownstreamStackBusLane[1][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane1_strm1_data          ( DownstreamStackBusLane[1][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane1_strm1_data_valid    ( DownstreamStackBusLane[1][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane2_strm0_ready         ( DownstreamStackBusLane[1][2].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane2_strm0_cntl          ( DownstreamStackBusLane[1][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane2_strm0_data          ( DownstreamStackBusLane[1][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane2_strm0_data_valid    ( DownstreamStackBusLane[1][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane2_strm1_ready         ( DownstreamStackBusLane[1][2].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane2_strm1_cntl          ( DownstreamStackBusLane[1][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane2_strm1_data          ( DownstreamStackBusLane[1][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane2_strm1_data_valid    ( DownstreamStackBusLane[1][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane3_strm0_ready         ( DownstreamStackBusLane[1][3].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane3_strm0_cntl          ( DownstreamStackBusLane[1][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane3_strm0_data          ( DownstreamStackBusLane[1][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane3_strm0_data_valid    ( DownstreamStackBusLane[1][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane3_strm1_ready         ( DownstreamStackBusLane[1][3].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane3_strm1_cntl          ( DownstreamStackBusLane[1][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane3_strm1_data          ( DownstreamStackBusLane[1][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane3_strm1_data_valid    ( DownstreamStackBusLane[1][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane4_strm0_ready         ( DownstreamStackBusLane[1][4].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane4_strm0_cntl          ( DownstreamStackBusLane[1][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane4_strm0_data          ( DownstreamStackBusLane[1][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane4_strm0_data_valid    ( DownstreamStackBusLane[1][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane4_strm1_ready         ( DownstreamStackBusLane[1][4].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane4_strm1_cntl          ( DownstreamStackBusLane[1][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane4_strm1_data          ( DownstreamStackBusLane[1][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane4_strm1_data_valid    ( DownstreamStackBusLane[1][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane5_strm0_ready         ( DownstreamStackBusLane[1][5].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane5_strm0_cntl          ( DownstreamStackBusLane[1][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane5_strm0_data          ( DownstreamStackBusLane[1][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane5_strm0_data_valid    ( DownstreamStackBusLane[1][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane5_strm1_ready         ( DownstreamStackBusLane[1][5].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane5_strm1_cntl          ( DownstreamStackBusLane[1][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane5_strm1_data          ( DownstreamStackBusLane[1][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane5_strm1_data_valid    ( DownstreamStackBusLane[1][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane6_strm0_ready         ( DownstreamStackBusLane[1][6].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane6_strm0_cntl          ( DownstreamStackBusLane[1][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane6_strm0_data          ( DownstreamStackBusLane[1][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane6_strm0_data_valid    ( DownstreamStackBusLane[1][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane6_strm1_ready         ( DownstreamStackBusLane[1][6].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane6_strm1_cntl          ( DownstreamStackBusLane[1][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane6_strm1_data          ( DownstreamStackBusLane[1][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane6_strm1_data_valid    ( DownstreamStackBusLane[1][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane7_strm0_ready         ( DownstreamStackBusLane[1][7].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane7_strm0_cntl          ( DownstreamStackBusLane[1][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane7_strm0_data          ( DownstreamStackBusLane[1][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane7_strm0_data_valid    ( DownstreamStackBusLane[1][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane7_strm1_ready         ( DownstreamStackBusLane[1][7].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane7_strm1_cntl          ( DownstreamStackBusLane[1][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane7_strm1_data          ( DownstreamStackBusLane[1][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane7_strm1_data_valid    ( DownstreamStackBusLane[1][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane8_strm0_ready         ( DownstreamStackBusLane[1][8].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane8_strm0_cntl          ( DownstreamStackBusLane[1][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane8_strm0_data          ( DownstreamStackBusLane[1][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane8_strm0_data_valid    ( DownstreamStackBusLane[1][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane8_strm1_ready         ( DownstreamStackBusLane[1][8].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane8_strm1_cntl          ( DownstreamStackBusLane[1][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane8_strm1_data          ( DownstreamStackBusLane[1][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane8_strm1_data_valid    ( DownstreamStackBusLane[1][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane9_strm0_ready         ( DownstreamStackBusLane[1][9].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane9_strm0_cntl          ( DownstreamStackBusLane[1][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane9_strm0_data          ( DownstreamStackBusLane[1][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane9_strm0_data_valid    ( DownstreamStackBusLane[1][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane9_strm1_ready         ( DownstreamStackBusLane[1][9].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane9_strm1_cntl          ( DownstreamStackBusLane[1][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane9_strm1_data          ( DownstreamStackBusLane[1][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane9_strm1_data_valid    ( DownstreamStackBusLane[1][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane10_strm0_ready         ( DownstreamStackBusLane[1][10].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane10_strm0_cntl          ( DownstreamStackBusLane[1][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane10_strm0_data          ( DownstreamStackBusLane[1][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane10_strm0_data_valid    ( DownstreamStackBusLane[1][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane10_strm1_ready         ( DownstreamStackBusLane[1][10].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane10_strm1_cntl          ( DownstreamStackBusLane[1][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane10_strm1_data          ( DownstreamStackBusLane[1][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane10_strm1_data_valid    ( DownstreamStackBusLane[1][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane11_strm0_ready         ( DownstreamStackBusLane[1][11].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane11_strm0_cntl          ( DownstreamStackBusLane[1][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane11_strm0_data          ( DownstreamStackBusLane[1][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane11_strm0_data_valid    ( DownstreamStackBusLane[1][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane11_strm1_ready         ( DownstreamStackBusLane[1][11].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane11_strm1_cntl          ( DownstreamStackBusLane[1][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane11_strm1_data          ( DownstreamStackBusLane[1][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane11_strm1_data_valid    ( DownstreamStackBusLane[1][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane12_strm0_ready         ( DownstreamStackBusLane[1][12].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane12_strm0_cntl          ( DownstreamStackBusLane[1][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane12_strm0_data          ( DownstreamStackBusLane[1][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane12_strm0_data_valid    ( DownstreamStackBusLane[1][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane12_strm1_ready         ( DownstreamStackBusLane[1][12].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane12_strm1_cntl          ( DownstreamStackBusLane[1][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane12_strm1_data          ( DownstreamStackBusLane[1][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane12_strm1_data_valid    ( DownstreamStackBusLane[1][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane13_strm0_ready         ( DownstreamStackBusLane[1][13].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane13_strm0_cntl          ( DownstreamStackBusLane[1][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane13_strm0_data          ( DownstreamStackBusLane[1][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane13_strm0_data_valid    ( DownstreamStackBusLane[1][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane13_strm1_ready         ( DownstreamStackBusLane[1][13].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane13_strm1_cntl          ( DownstreamStackBusLane[1][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane13_strm1_data          ( DownstreamStackBusLane[1][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane13_strm1_data_valid    ( DownstreamStackBusLane[1][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane14_strm0_ready         ( DownstreamStackBusLane[1][14].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane14_strm0_cntl          ( DownstreamStackBusLane[1][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane14_strm0_data          ( DownstreamStackBusLane[1][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane14_strm0_data_valid    ( DownstreamStackBusLane[1][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane14_strm1_ready         ( DownstreamStackBusLane[1][14].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane14_strm1_cntl          ( DownstreamStackBusLane[1][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane14_strm1_data          ( DownstreamStackBusLane[1][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane14_strm1_data_valid    ( DownstreamStackBusLane[1][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane15_strm0_ready         ( DownstreamStackBusLane[1][15].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane15_strm0_cntl          ( DownstreamStackBusLane[1][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane15_strm0_data          ( DownstreamStackBusLane[1][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane15_strm0_data_valid    ( DownstreamStackBusLane[1][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane15_strm1_ready         ( DownstreamStackBusLane[1][15].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane15_strm1_cntl          ( DownstreamStackBusLane[1][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane15_strm1_data          ( DownstreamStackBusLane[1][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane15_strm1_data_valid    ( DownstreamStackBusLane[1][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane16_strm0_ready         ( DownstreamStackBusLane[1][16].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane16_strm0_cntl          ( DownstreamStackBusLane[1][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane16_strm0_data          ( DownstreamStackBusLane[1][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane16_strm0_data_valid    ( DownstreamStackBusLane[1][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane16_strm1_ready         ( DownstreamStackBusLane[1][16].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane16_strm1_cntl          ( DownstreamStackBusLane[1][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane16_strm1_data          ( DownstreamStackBusLane[1][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane16_strm1_data_valid    ( DownstreamStackBusLane[1][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane17_strm0_ready         ( DownstreamStackBusLane[1][17].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane17_strm0_cntl          ( DownstreamStackBusLane[1][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane17_strm0_data          ( DownstreamStackBusLane[1][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane17_strm0_data_valid    ( DownstreamStackBusLane[1][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane17_strm1_ready         ( DownstreamStackBusLane[1][17].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane17_strm1_cntl          ( DownstreamStackBusLane[1][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane17_strm1_data          ( DownstreamStackBusLane[1][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane17_strm1_data_valid    ( DownstreamStackBusLane[1][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane18_strm0_ready         ( DownstreamStackBusLane[1][18].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane18_strm0_cntl          ( DownstreamStackBusLane[1][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane18_strm0_data          ( DownstreamStackBusLane[1][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane18_strm0_data_valid    ( DownstreamStackBusLane[1][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane18_strm1_ready         ( DownstreamStackBusLane[1][18].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane18_strm1_cntl          ( DownstreamStackBusLane[1][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane18_strm1_data          ( DownstreamStackBusLane[1][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane18_strm1_data_valid    ( DownstreamStackBusLane[1][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane19_strm0_ready         ( DownstreamStackBusLane[1][19].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane19_strm0_cntl          ( DownstreamStackBusLane[1][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane19_strm0_data          ( DownstreamStackBusLane[1][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane19_strm0_data_valid    ( DownstreamStackBusLane[1][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane19_strm1_ready         ( DownstreamStackBusLane[1][19].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane19_strm1_cntl          ( DownstreamStackBusLane[1][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane19_strm1_data          ( DownstreamStackBusLane[1][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane19_strm1_data_valid    ( DownstreamStackBusLane[1][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane20_strm0_ready         ( DownstreamStackBusLane[1][20].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane20_strm0_cntl          ( DownstreamStackBusLane[1][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane20_strm0_data          ( DownstreamStackBusLane[1][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane20_strm0_data_valid    ( DownstreamStackBusLane[1][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane20_strm1_ready         ( DownstreamStackBusLane[1][20].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane20_strm1_cntl          ( DownstreamStackBusLane[1][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane20_strm1_data          ( DownstreamStackBusLane[1][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane20_strm1_data_valid    ( DownstreamStackBusLane[1][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane21_strm0_ready         ( DownstreamStackBusLane[1][21].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane21_strm0_cntl          ( DownstreamStackBusLane[1][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane21_strm0_data          ( DownstreamStackBusLane[1][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane21_strm0_data_valid    ( DownstreamStackBusLane[1][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane21_strm1_ready         ( DownstreamStackBusLane[1][21].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane21_strm1_cntl          ( DownstreamStackBusLane[1][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane21_strm1_data          ( DownstreamStackBusLane[1][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane21_strm1_data_valid    ( DownstreamStackBusLane[1][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane22_strm0_ready         ( DownstreamStackBusLane[1][22].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane22_strm0_cntl          ( DownstreamStackBusLane[1][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane22_strm0_data          ( DownstreamStackBusLane[1][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane22_strm0_data_valid    ( DownstreamStackBusLane[1][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane22_strm1_ready         ( DownstreamStackBusLane[1][22].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane22_strm1_cntl          ( DownstreamStackBusLane[1][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane22_strm1_data          ( DownstreamStackBusLane[1][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane22_strm1_data_valid    ( DownstreamStackBusLane[1][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane23_strm0_ready         ( DownstreamStackBusLane[1][23].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane23_strm0_cntl          ( DownstreamStackBusLane[1][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane23_strm0_data          ( DownstreamStackBusLane[1][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane23_strm0_data_valid    ( DownstreamStackBusLane[1][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane23_strm1_ready         ( DownstreamStackBusLane[1][23].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane23_strm1_cntl          ( DownstreamStackBusLane[1][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane23_strm1_data          ( DownstreamStackBusLane[1][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane23_strm1_data_valid    ( DownstreamStackBusLane[1][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane24_strm0_ready         ( DownstreamStackBusLane[1][24].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane24_strm0_cntl          ( DownstreamStackBusLane[1][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane24_strm0_data          ( DownstreamStackBusLane[1][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane24_strm0_data_valid    ( DownstreamStackBusLane[1][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane24_strm1_ready         ( DownstreamStackBusLane[1][24].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane24_strm1_cntl          ( DownstreamStackBusLane[1][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane24_strm1_data          ( DownstreamStackBusLane[1][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane24_strm1_data_valid    ( DownstreamStackBusLane[1][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane25_strm0_ready         ( DownstreamStackBusLane[1][25].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane25_strm0_cntl          ( DownstreamStackBusLane[1][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane25_strm0_data          ( DownstreamStackBusLane[1][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane25_strm0_data_valid    ( DownstreamStackBusLane[1][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane25_strm1_ready         ( DownstreamStackBusLane[1][25].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane25_strm1_cntl          ( DownstreamStackBusLane[1][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane25_strm1_data          ( DownstreamStackBusLane[1][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane25_strm1_data_valid    ( DownstreamStackBusLane[1][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane26_strm0_ready         ( DownstreamStackBusLane[1][26].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane26_strm0_cntl          ( DownstreamStackBusLane[1][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane26_strm0_data          ( DownstreamStackBusLane[1][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane26_strm0_data_valid    ( DownstreamStackBusLane[1][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane26_strm1_ready         ( DownstreamStackBusLane[1][26].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane26_strm1_cntl          ( DownstreamStackBusLane[1][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane26_strm1_data          ( DownstreamStackBusLane[1][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane26_strm1_data_valid    ( DownstreamStackBusLane[1][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane27_strm0_ready         ( DownstreamStackBusLane[1][27].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane27_strm0_cntl          ( DownstreamStackBusLane[1][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane27_strm0_data          ( DownstreamStackBusLane[1][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane27_strm0_data_valid    ( DownstreamStackBusLane[1][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane27_strm1_ready         ( DownstreamStackBusLane[1][27].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane27_strm1_cntl          ( DownstreamStackBusLane[1][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane27_strm1_data          ( DownstreamStackBusLane[1][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane27_strm1_data_valid    ( DownstreamStackBusLane[1][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane28_strm0_ready         ( DownstreamStackBusLane[1][28].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane28_strm0_cntl          ( DownstreamStackBusLane[1][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane28_strm0_data          ( DownstreamStackBusLane[1][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane28_strm0_data_valid    ( DownstreamStackBusLane[1][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane28_strm1_ready         ( DownstreamStackBusLane[1][28].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane28_strm1_cntl          ( DownstreamStackBusLane[1][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane28_strm1_data          ( DownstreamStackBusLane[1][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane28_strm1_data_valid    ( DownstreamStackBusLane[1][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane29_strm0_ready         ( DownstreamStackBusLane[1][29].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane29_strm0_cntl          ( DownstreamStackBusLane[1][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane29_strm0_data          ( DownstreamStackBusLane[1][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane29_strm0_data_valid    ( DownstreamStackBusLane[1][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane29_strm1_ready         ( DownstreamStackBusLane[1][29].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane29_strm1_cntl          ( DownstreamStackBusLane[1][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane29_strm1_data          ( DownstreamStackBusLane[1][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane29_strm1_data_valid    ( DownstreamStackBusLane[1][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane30_strm0_ready         ( DownstreamStackBusLane[1][30].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane30_strm0_cntl          ( DownstreamStackBusLane[1][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane30_strm0_data          ( DownstreamStackBusLane[1][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane30_strm0_data_valid    ( DownstreamStackBusLane[1][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane30_strm1_ready         ( DownstreamStackBusLane[1][30].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane30_strm1_cntl          ( DownstreamStackBusLane[1][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane30_strm1_data          ( DownstreamStackBusLane[1][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane30_strm1_data_valid    ( DownstreamStackBusLane[1][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane31_strm0_ready         ( DownstreamStackBusLane[1][31].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane31_strm0_cntl          ( DownstreamStackBusLane[1][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane31_strm0_data          ( DownstreamStackBusLane[1][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane31_strm0_data_valid    ( DownstreamStackBusLane[1][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane31_strm1_ready         ( DownstreamStackBusLane[1][31].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane31_strm1_cntl          ( DownstreamStackBusLane[1][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane31_strm1_data          ( DownstreamStackBusLane[1][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane31_strm1_data_valid    ( DownstreamStackBusLane[1][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane0_strm0_ready         ( DownstreamStackBusLane[2][0].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane0_strm0_cntl          ( DownstreamStackBusLane[2][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane0_strm0_data          ( DownstreamStackBusLane[2][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane0_strm0_data_valid    ( DownstreamStackBusLane[2][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane0_strm1_ready         ( DownstreamStackBusLane[2][0].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane0_strm1_cntl          ( DownstreamStackBusLane[2][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane0_strm1_data          ( DownstreamStackBusLane[2][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane0_strm1_data_valid    ( DownstreamStackBusLane[2][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane1_strm0_ready         ( DownstreamStackBusLane[2][1].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane1_strm0_cntl          ( DownstreamStackBusLane[2][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane1_strm0_data          ( DownstreamStackBusLane[2][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane1_strm0_data_valid    ( DownstreamStackBusLane[2][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane1_strm1_ready         ( DownstreamStackBusLane[2][1].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane1_strm1_cntl          ( DownstreamStackBusLane[2][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane1_strm1_data          ( DownstreamStackBusLane[2][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane1_strm1_data_valid    ( DownstreamStackBusLane[2][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane2_strm0_ready         ( DownstreamStackBusLane[2][2].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane2_strm0_cntl          ( DownstreamStackBusLane[2][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane2_strm0_data          ( DownstreamStackBusLane[2][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane2_strm0_data_valid    ( DownstreamStackBusLane[2][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane2_strm1_ready         ( DownstreamStackBusLane[2][2].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane2_strm1_cntl          ( DownstreamStackBusLane[2][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane2_strm1_data          ( DownstreamStackBusLane[2][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane2_strm1_data_valid    ( DownstreamStackBusLane[2][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane3_strm0_ready         ( DownstreamStackBusLane[2][3].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane3_strm0_cntl          ( DownstreamStackBusLane[2][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane3_strm0_data          ( DownstreamStackBusLane[2][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane3_strm0_data_valid    ( DownstreamStackBusLane[2][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane3_strm1_ready         ( DownstreamStackBusLane[2][3].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane3_strm1_cntl          ( DownstreamStackBusLane[2][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane3_strm1_data          ( DownstreamStackBusLane[2][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane3_strm1_data_valid    ( DownstreamStackBusLane[2][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane4_strm0_ready         ( DownstreamStackBusLane[2][4].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane4_strm0_cntl          ( DownstreamStackBusLane[2][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane4_strm0_data          ( DownstreamStackBusLane[2][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane4_strm0_data_valid    ( DownstreamStackBusLane[2][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane4_strm1_ready         ( DownstreamStackBusLane[2][4].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane4_strm1_cntl          ( DownstreamStackBusLane[2][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane4_strm1_data          ( DownstreamStackBusLane[2][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane4_strm1_data_valid    ( DownstreamStackBusLane[2][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane5_strm0_ready         ( DownstreamStackBusLane[2][5].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane5_strm0_cntl          ( DownstreamStackBusLane[2][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane5_strm0_data          ( DownstreamStackBusLane[2][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane5_strm0_data_valid    ( DownstreamStackBusLane[2][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane5_strm1_ready         ( DownstreamStackBusLane[2][5].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane5_strm1_cntl          ( DownstreamStackBusLane[2][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane5_strm1_data          ( DownstreamStackBusLane[2][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane5_strm1_data_valid    ( DownstreamStackBusLane[2][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane6_strm0_ready         ( DownstreamStackBusLane[2][6].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane6_strm0_cntl          ( DownstreamStackBusLane[2][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane6_strm0_data          ( DownstreamStackBusLane[2][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane6_strm0_data_valid    ( DownstreamStackBusLane[2][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane6_strm1_ready         ( DownstreamStackBusLane[2][6].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane6_strm1_cntl          ( DownstreamStackBusLane[2][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane6_strm1_data          ( DownstreamStackBusLane[2][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane6_strm1_data_valid    ( DownstreamStackBusLane[2][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane7_strm0_ready         ( DownstreamStackBusLane[2][7].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane7_strm0_cntl          ( DownstreamStackBusLane[2][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane7_strm0_data          ( DownstreamStackBusLane[2][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane7_strm0_data_valid    ( DownstreamStackBusLane[2][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane7_strm1_ready         ( DownstreamStackBusLane[2][7].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane7_strm1_cntl          ( DownstreamStackBusLane[2][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane7_strm1_data          ( DownstreamStackBusLane[2][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane7_strm1_data_valid    ( DownstreamStackBusLane[2][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane8_strm0_ready         ( DownstreamStackBusLane[2][8].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane8_strm0_cntl          ( DownstreamStackBusLane[2][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane8_strm0_data          ( DownstreamStackBusLane[2][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane8_strm0_data_valid    ( DownstreamStackBusLane[2][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane8_strm1_ready         ( DownstreamStackBusLane[2][8].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane8_strm1_cntl          ( DownstreamStackBusLane[2][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane8_strm1_data          ( DownstreamStackBusLane[2][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane8_strm1_data_valid    ( DownstreamStackBusLane[2][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane9_strm0_ready         ( DownstreamStackBusLane[2][9].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane9_strm0_cntl          ( DownstreamStackBusLane[2][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane9_strm0_data          ( DownstreamStackBusLane[2][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane9_strm0_data_valid    ( DownstreamStackBusLane[2][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane9_strm1_ready         ( DownstreamStackBusLane[2][9].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane9_strm1_cntl          ( DownstreamStackBusLane[2][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane9_strm1_data          ( DownstreamStackBusLane[2][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane9_strm1_data_valid    ( DownstreamStackBusLane[2][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane10_strm0_ready         ( DownstreamStackBusLane[2][10].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane10_strm0_cntl          ( DownstreamStackBusLane[2][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane10_strm0_data          ( DownstreamStackBusLane[2][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane10_strm0_data_valid    ( DownstreamStackBusLane[2][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane10_strm1_ready         ( DownstreamStackBusLane[2][10].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane10_strm1_cntl          ( DownstreamStackBusLane[2][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane10_strm1_data          ( DownstreamStackBusLane[2][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane10_strm1_data_valid    ( DownstreamStackBusLane[2][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane11_strm0_ready         ( DownstreamStackBusLane[2][11].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane11_strm0_cntl          ( DownstreamStackBusLane[2][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane11_strm0_data          ( DownstreamStackBusLane[2][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane11_strm0_data_valid    ( DownstreamStackBusLane[2][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane11_strm1_ready         ( DownstreamStackBusLane[2][11].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane11_strm1_cntl          ( DownstreamStackBusLane[2][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane11_strm1_data          ( DownstreamStackBusLane[2][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane11_strm1_data_valid    ( DownstreamStackBusLane[2][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane12_strm0_ready         ( DownstreamStackBusLane[2][12].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane12_strm0_cntl          ( DownstreamStackBusLane[2][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane12_strm0_data          ( DownstreamStackBusLane[2][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane12_strm0_data_valid    ( DownstreamStackBusLane[2][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane12_strm1_ready         ( DownstreamStackBusLane[2][12].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane12_strm1_cntl          ( DownstreamStackBusLane[2][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane12_strm1_data          ( DownstreamStackBusLane[2][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane12_strm1_data_valid    ( DownstreamStackBusLane[2][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane13_strm0_ready         ( DownstreamStackBusLane[2][13].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane13_strm0_cntl          ( DownstreamStackBusLane[2][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane13_strm0_data          ( DownstreamStackBusLane[2][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane13_strm0_data_valid    ( DownstreamStackBusLane[2][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane13_strm1_ready         ( DownstreamStackBusLane[2][13].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane13_strm1_cntl          ( DownstreamStackBusLane[2][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane13_strm1_data          ( DownstreamStackBusLane[2][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane13_strm1_data_valid    ( DownstreamStackBusLane[2][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane14_strm0_ready         ( DownstreamStackBusLane[2][14].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane14_strm0_cntl          ( DownstreamStackBusLane[2][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane14_strm0_data          ( DownstreamStackBusLane[2][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane14_strm0_data_valid    ( DownstreamStackBusLane[2][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane14_strm1_ready         ( DownstreamStackBusLane[2][14].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane14_strm1_cntl          ( DownstreamStackBusLane[2][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane14_strm1_data          ( DownstreamStackBusLane[2][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane14_strm1_data_valid    ( DownstreamStackBusLane[2][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane15_strm0_ready         ( DownstreamStackBusLane[2][15].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane15_strm0_cntl          ( DownstreamStackBusLane[2][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane15_strm0_data          ( DownstreamStackBusLane[2][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane15_strm0_data_valid    ( DownstreamStackBusLane[2][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane15_strm1_ready         ( DownstreamStackBusLane[2][15].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane15_strm1_cntl          ( DownstreamStackBusLane[2][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane15_strm1_data          ( DownstreamStackBusLane[2][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane15_strm1_data_valid    ( DownstreamStackBusLane[2][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane16_strm0_ready         ( DownstreamStackBusLane[2][16].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane16_strm0_cntl          ( DownstreamStackBusLane[2][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane16_strm0_data          ( DownstreamStackBusLane[2][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane16_strm0_data_valid    ( DownstreamStackBusLane[2][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane16_strm1_ready         ( DownstreamStackBusLane[2][16].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane16_strm1_cntl          ( DownstreamStackBusLane[2][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane16_strm1_data          ( DownstreamStackBusLane[2][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane16_strm1_data_valid    ( DownstreamStackBusLane[2][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane17_strm0_ready         ( DownstreamStackBusLane[2][17].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane17_strm0_cntl          ( DownstreamStackBusLane[2][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane17_strm0_data          ( DownstreamStackBusLane[2][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane17_strm0_data_valid    ( DownstreamStackBusLane[2][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane17_strm1_ready         ( DownstreamStackBusLane[2][17].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane17_strm1_cntl          ( DownstreamStackBusLane[2][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane17_strm1_data          ( DownstreamStackBusLane[2][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane17_strm1_data_valid    ( DownstreamStackBusLane[2][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane18_strm0_ready         ( DownstreamStackBusLane[2][18].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane18_strm0_cntl          ( DownstreamStackBusLane[2][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane18_strm0_data          ( DownstreamStackBusLane[2][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane18_strm0_data_valid    ( DownstreamStackBusLane[2][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane18_strm1_ready         ( DownstreamStackBusLane[2][18].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane18_strm1_cntl          ( DownstreamStackBusLane[2][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane18_strm1_data          ( DownstreamStackBusLane[2][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane18_strm1_data_valid    ( DownstreamStackBusLane[2][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane19_strm0_ready         ( DownstreamStackBusLane[2][19].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane19_strm0_cntl          ( DownstreamStackBusLane[2][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane19_strm0_data          ( DownstreamStackBusLane[2][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane19_strm0_data_valid    ( DownstreamStackBusLane[2][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane19_strm1_ready         ( DownstreamStackBusLane[2][19].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane19_strm1_cntl          ( DownstreamStackBusLane[2][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane19_strm1_data          ( DownstreamStackBusLane[2][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane19_strm1_data_valid    ( DownstreamStackBusLane[2][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane20_strm0_ready         ( DownstreamStackBusLane[2][20].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane20_strm0_cntl          ( DownstreamStackBusLane[2][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane20_strm0_data          ( DownstreamStackBusLane[2][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane20_strm0_data_valid    ( DownstreamStackBusLane[2][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane20_strm1_ready         ( DownstreamStackBusLane[2][20].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane20_strm1_cntl          ( DownstreamStackBusLane[2][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane20_strm1_data          ( DownstreamStackBusLane[2][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane20_strm1_data_valid    ( DownstreamStackBusLane[2][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane21_strm0_ready         ( DownstreamStackBusLane[2][21].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane21_strm0_cntl          ( DownstreamStackBusLane[2][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane21_strm0_data          ( DownstreamStackBusLane[2][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane21_strm0_data_valid    ( DownstreamStackBusLane[2][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane21_strm1_ready         ( DownstreamStackBusLane[2][21].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane21_strm1_cntl          ( DownstreamStackBusLane[2][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane21_strm1_data          ( DownstreamStackBusLane[2][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane21_strm1_data_valid    ( DownstreamStackBusLane[2][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane22_strm0_ready         ( DownstreamStackBusLane[2][22].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane22_strm0_cntl          ( DownstreamStackBusLane[2][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane22_strm0_data          ( DownstreamStackBusLane[2][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane22_strm0_data_valid    ( DownstreamStackBusLane[2][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane22_strm1_ready         ( DownstreamStackBusLane[2][22].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane22_strm1_cntl          ( DownstreamStackBusLane[2][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane22_strm1_data          ( DownstreamStackBusLane[2][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane22_strm1_data_valid    ( DownstreamStackBusLane[2][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane23_strm0_ready         ( DownstreamStackBusLane[2][23].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane23_strm0_cntl          ( DownstreamStackBusLane[2][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane23_strm0_data          ( DownstreamStackBusLane[2][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane23_strm0_data_valid    ( DownstreamStackBusLane[2][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane23_strm1_ready         ( DownstreamStackBusLane[2][23].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane23_strm1_cntl          ( DownstreamStackBusLane[2][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane23_strm1_data          ( DownstreamStackBusLane[2][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane23_strm1_data_valid    ( DownstreamStackBusLane[2][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane24_strm0_ready         ( DownstreamStackBusLane[2][24].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane24_strm0_cntl          ( DownstreamStackBusLane[2][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane24_strm0_data          ( DownstreamStackBusLane[2][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane24_strm0_data_valid    ( DownstreamStackBusLane[2][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane24_strm1_ready         ( DownstreamStackBusLane[2][24].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane24_strm1_cntl          ( DownstreamStackBusLane[2][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane24_strm1_data          ( DownstreamStackBusLane[2][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane24_strm1_data_valid    ( DownstreamStackBusLane[2][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane25_strm0_ready         ( DownstreamStackBusLane[2][25].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane25_strm0_cntl          ( DownstreamStackBusLane[2][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane25_strm0_data          ( DownstreamStackBusLane[2][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane25_strm0_data_valid    ( DownstreamStackBusLane[2][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane25_strm1_ready         ( DownstreamStackBusLane[2][25].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane25_strm1_cntl          ( DownstreamStackBusLane[2][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane25_strm1_data          ( DownstreamStackBusLane[2][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane25_strm1_data_valid    ( DownstreamStackBusLane[2][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane26_strm0_ready         ( DownstreamStackBusLane[2][26].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane26_strm0_cntl          ( DownstreamStackBusLane[2][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane26_strm0_data          ( DownstreamStackBusLane[2][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane26_strm0_data_valid    ( DownstreamStackBusLane[2][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane26_strm1_ready         ( DownstreamStackBusLane[2][26].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane26_strm1_cntl          ( DownstreamStackBusLane[2][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane26_strm1_data          ( DownstreamStackBusLane[2][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane26_strm1_data_valid    ( DownstreamStackBusLane[2][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane27_strm0_ready         ( DownstreamStackBusLane[2][27].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane27_strm0_cntl          ( DownstreamStackBusLane[2][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane27_strm0_data          ( DownstreamStackBusLane[2][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane27_strm0_data_valid    ( DownstreamStackBusLane[2][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane27_strm1_ready         ( DownstreamStackBusLane[2][27].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane27_strm1_cntl          ( DownstreamStackBusLane[2][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane27_strm1_data          ( DownstreamStackBusLane[2][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane27_strm1_data_valid    ( DownstreamStackBusLane[2][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane28_strm0_ready         ( DownstreamStackBusLane[2][28].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane28_strm0_cntl          ( DownstreamStackBusLane[2][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane28_strm0_data          ( DownstreamStackBusLane[2][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane28_strm0_data_valid    ( DownstreamStackBusLane[2][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane28_strm1_ready         ( DownstreamStackBusLane[2][28].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane28_strm1_cntl          ( DownstreamStackBusLane[2][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane28_strm1_data          ( DownstreamStackBusLane[2][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane28_strm1_data_valid    ( DownstreamStackBusLane[2][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane29_strm0_ready         ( DownstreamStackBusLane[2][29].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane29_strm0_cntl          ( DownstreamStackBusLane[2][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane29_strm0_data          ( DownstreamStackBusLane[2][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane29_strm0_data_valid    ( DownstreamStackBusLane[2][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane29_strm1_ready         ( DownstreamStackBusLane[2][29].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane29_strm1_cntl          ( DownstreamStackBusLane[2][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane29_strm1_data          ( DownstreamStackBusLane[2][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane29_strm1_data_valid    ( DownstreamStackBusLane[2][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane30_strm0_ready         ( DownstreamStackBusLane[2][30].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane30_strm0_cntl          ( DownstreamStackBusLane[2][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane30_strm0_data          ( DownstreamStackBusLane[2][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane30_strm0_data_valid    ( DownstreamStackBusLane[2][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane30_strm1_ready         ( DownstreamStackBusLane[2][30].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane30_strm1_cntl          ( DownstreamStackBusLane[2][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane30_strm1_data          ( DownstreamStackBusLane[2][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane30_strm1_data_valid    ( DownstreamStackBusLane[2][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane31_strm0_ready         ( DownstreamStackBusLane[2][31].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane31_strm0_cntl          ( DownstreamStackBusLane[2][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane31_strm0_data          ( DownstreamStackBusLane[2][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane31_strm0_data_valid    ( DownstreamStackBusLane[2][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane31_strm1_ready         ( DownstreamStackBusLane[2][31].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane31_strm1_cntl          ( DownstreamStackBusLane[2][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane31_strm1_data          ( DownstreamStackBusLane[2][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane31_strm1_data_valid    ( DownstreamStackBusLane[2][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane0_strm0_ready         ( DownstreamStackBusLane[3][0].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane0_strm0_cntl          ( DownstreamStackBusLane[3][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane0_strm0_data          ( DownstreamStackBusLane[3][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane0_strm0_data_valid    ( DownstreamStackBusLane[3][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane0_strm1_ready         ( DownstreamStackBusLane[3][0].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane0_strm1_cntl          ( DownstreamStackBusLane[3][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane0_strm1_data          ( DownstreamStackBusLane[3][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane0_strm1_data_valid    ( DownstreamStackBusLane[3][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane1_strm0_ready         ( DownstreamStackBusLane[3][1].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane1_strm0_cntl          ( DownstreamStackBusLane[3][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane1_strm0_data          ( DownstreamStackBusLane[3][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane1_strm0_data_valid    ( DownstreamStackBusLane[3][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane1_strm1_ready         ( DownstreamStackBusLane[3][1].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane1_strm1_cntl          ( DownstreamStackBusLane[3][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane1_strm1_data          ( DownstreamStackBusLane[3][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane1_strm1_data_valid    ( DownstreamStackBusLane[3][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane2_strm0_ready         ( DownstreamStackBusLane[3][2].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane2_strm0_cntl          ( DownstreamStackBusLane[3][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane2_strm0_data          ( DownstreamStackBusLane[3][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane2_strm0_data_valid    ( DownstreamStackBusLane[3][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane2_strm1_ready         ( DownstreamStackBusLane[3][2].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane2_strm1_cntl          ( DownstreamStackBusLane[3][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane2_strm1_data          ( DownstreamStackBusLane[3][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane2_strm1_data_valid    ( DownstreamStackBusLane[3][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane3_strm0_ready         ( DownstreamStackBusLane[3][3].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane3_strm0_cntl          ( DownstreamStackBusLane[3][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane3_strm0_data          ( DownstreamStackBusLane[3][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane3_strm0_data_valid    ( DownstreamStackBusLane[3][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane3_strm1_ready         ( DownstreamStackBusLane[3][3].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane3_strm1_cntl          ( DownstreamStackBusLane[3][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane3_strm1_data          ( DownstreamStackBusLane[3][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane3_strm1_data_valid    ( DownstreamStackBusLane[3][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane4_strm0_ready         ( DownstreamStackBusLane[3][4].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane4_strm0_cntl          ( DownstreamStackBusLane[3][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane4_strm0_data          ( DownstreamStackBusLane[3][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane4_strm0_data_valid    ( DownstreamStackBusLane[3][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane4_strm1_ready         ( DownstreamStackBusLane[3][4].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane4_strm1_cntl          ( DownstreamStackBusLane[3][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane4_strm1_data          ( DownstreamStackBusLane[3][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane4_strm1_data_valid    ( DownstreamStackBusLane[3][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane5_strm0_ready         ( DownstreamStackBusLane[3][5].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane5_strm0_cntl          ( DownstreamStackBusLane[3][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane5_strm0_data          ( DownstreamStackBusLane[3][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane5_strm0_data_valid    ( DownstreamStackBusLane[3][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane5_strm1_ready         ( DownstreamStackBusLane[3][5].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane5_strm1_cntl          ( DownstreamStackBusLane[3][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane5_strm1_data          ( DownstreamStackBusLane[3][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane5_strm1_data_valid    ( DownstreamStackBusLane[3][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane6_strm0_ready         ( DownstreamStackBusLane[3][6].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane6_strm0_cntl          ( DownstreamStackBusLane[3][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane6_strm0_data          ( DownstreamStackBusLane[3][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane6_strm0_data_valid    ( DownstreamStackBusLane[3][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane6_strm1_ready         ( DownstreamStackBusLane[3][6].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane6_strm1_cntl          ( DownstreamStackBusLane[3][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane6_strm1_data          ( DownstreamStackBusLane[3][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane6_strm1_data_valid    ( DownstreamStackBusLane[3][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane7_strm0_ready         ( DownstreamStackBusLane[3][7].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane7_strm0_cntl          ( DownstreamStackBusLane[3][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane7_strm0_data          ( DownstreamStackBusLane[3][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane7_strm0_data_valid    ( DownstreamStackBusLane[3][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane7_strm1_ready         ( DownstreamStackBusLane[3][7].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane7_strm1_cntl          ( DownstreamStackBusLane[3][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane7_strm1_data          ( DownstreamStackBusLane[3][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane7_strm1_data_valid    ( DownstreamStackBusLane[3][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane8_strm0_ready         ( DownstreamStackBusLane[3][8].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane8_strm0_cntl          ( DownstreamStackBusLane[3][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane8_strm0_data          ( DownstreamStackBusLane[3][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane8_strm0_data_valid    ( DownstreamStackBusLane[3][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane8_strm1_ready         ( DownstreamStackBusLane[3][8].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane8_strm1_cntl          ( DownstreamStackBusLane[3][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane8_strm1_data          ( DownstreamStackBusLane[3][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane8_strm1_data_valid    ( DownstreamStackBusLane[3][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane9_strm0_ready         ( DownstreamStackBusLane[3][9].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane9_strm0_cntl          ( DownstreamStackBusLane[3][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane9_strm0_data          ( DownstreamStackBusLane[3][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane9_strm0_data_valid    ( DownstreamStackBusLane[3][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane9_strm1_ready         ( DownstreamStackBusLane[3][9].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane9_strm1_cntl          ( DownstreamStackBusLane[3][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane9_strm1_data          ( DownstreamStackBusLane[3][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane9_strm1_data_valid    ( DownstreamStackBusLane[3][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane10_strm0_ready         ( DownstreamStackBusLane[3][10].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane10_strm0_cntl          ( DownstreamStackBusLane[3][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane10_strm0_data          ( DownstreamStackBusLane[3][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane10_strm0_data_valid    ( DownstreamStackBusLane[3][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane10_strm1_ready         ( DownstreamStackBusLane[3][10].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane10_strm1_cntl          ( DownstreamStackBusLane[3][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane10_strm1_data          ( DownstreamStackBusLane[3][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane10_strm1_data_valid    ( DownstreamStackBusLane[3][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane11_strm0_ready         ( DownstreamStackBusLane[3][11].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane11_strm0_cntl          ( DownstreamStackBusLane[3][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane11_strm0_data          ( DownstreamStackBusLane[3][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane11_strm0_data_valid    ( DownstreamStackBusLane[3][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane11_strm1_ready         ( DownstreamStackBusLane[3][11].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane11_strm1_cntl          ( DownstreamStackBusLane[3][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane11_strm1_data          ( DownstreamStackBusLane[3][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane11_strm1_data_valid    ( DownstreamStackBusLane[3][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane12_strm0_ready         ( DownstreamStackBusLane[3][12].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane12_strm0_cntl          ( DownstreamStackBusLane[3][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane12_strm0_data          ( DownstreamStackBusLane[3][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane12_strm0_data_valid    ( DownstreamStackBusLane[3][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane12_strm1_ready         ( DownstreamStackBusLane[3][12].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane12_strm1_cntl          ( DownstreamStackBusLane[3][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane12_strm1_data          ( DownstreamStackBusLane[3][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane12_strm1_data_valid    ( DownstreamStackBusLane[3][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane13_strm0_ready         ( DownstreamStackBusLane[3][13].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane13_strm0_cntl          ( DownstreamStackBusLane[3][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane13_strm0_data          ( DownstreamStackBusLane[3][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane13_strm0_data_valid    ( DownstreamStackBusLane[3][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane13_strm1_ready         ( DownstreamStackBusLane[3][13].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane13_strm1_cntl          ( DownstreamStackBusLane[3][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane13_strm1_data          ( DownstreamStackBusLane[3][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane13_strm1_data_valid    ( DownstreamStackBusLane[3][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane14_strm0_ready         ( DownstreamStackBusLane[3][14].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane14_strm0_cntl          ( DownstreamStackBusLane[3][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane14_strm0_data          ( DownstreamStackBusLane[3][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane14_strm0_data_valid    ( DownstreamStackBusLane[3][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane14_strm1_ready         ( DownstreamStackBusLane[3][14].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane14_strm1_cntl          ( DownstreamStackBusLane[3][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane14_strm1_data          ( DownstreamStackBusLane[3][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane14_strm1_data_valid    ( DownstreamStackBusLane[3][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane15_strm0_ready         ( DownstreamStackBusLane[3][15].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane15_strm0_cntl          ( DownstreamStackBusLane[3][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane15_strm0_data          ( DownstreamStackBusLane[3][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane15_strm0_data_valid    ( DownstreamStackBusLane[3][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane15_strm1_ready         ( DownstreamStackBusLane[3][15].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane15_strm1_cntl          ( DownstreamStackBusLane[3][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane15_strm1_data          ( DownstreamStackBusLane[3][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane15_strm1_data_valid    ( DownstreamStackBusLane[3][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane16_strm0_ready         ( DownstreamStackBusLane[3][16].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane16_strm0_cntl          ( DownstreamStackBusLane[3][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane16_strm0_data          ( DownstreamStackBusLane[3][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane16_strm0_data_valid    ( DownstreamStackBusLane[3][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane16_strm1_ready         ( DownstreamStackBusLane[3][16].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane16_strm1_cntl          ( DownstreamStackBusLane[3][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane16_strm1_data          ( DownstreamStackBusLane[3][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane16_strm1_data_valid    ( DownstreamStackBusLane[3][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane17_strm0_ready         ( DownstreamStackBusLane[3][17].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane17_strm0_cntl          ( DownstreamStackBusLane[3][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane17_strm0_data          ( DownstreamStackBusLane[3][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane17_strm0_data_valid    ( DownstreamStackBusLane[3][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane17_strm1_ready         ( DownstreamStackBusLane[3][17].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane17_strm1_cntl          ( DownstreamStackBusLane[3][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane17_strm1_data          ( DownstreamStackBusLane[3][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane17_strm1_data_valid    ( DownstreamStackBusLane[3][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane18_strm0_ready         ( DownstreamStackBusLane[3][18].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane18_strm0_cntl          ( DownstreamStackBusLane[3][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane18_strm0_data          ( DownstreamStackBusLane[3][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane18_strm0_data_valid    ( DownstreamStackBusLane[3][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane18_strm1_ready         ( DownstreamStackBusLane[3][18].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane18_strm1_cntl          ( DownstreamStackBusLane[3][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane18_strm1_data          ( DownstreamStackBusLane[3][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane18_strm1_data_valid    ( DownstreamStackBusLane[3][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane19_strm0_ready         ( DownstreamStackBusLane[3][19].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane19_strm0_cntl          ( DownstreamStackBusLane[3][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane19_strm0_data          ( DownstreamStackBusLane[3][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane19_strm0_data_valid    ( DownstreamStackBusLane[3][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane19_strm1_ready         ( DownstreamStackBusLane[3][19].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane19_strm1_cntl          ( DownstreamStackBusLane[3][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane19_strm1_data          ( DownstreamStackBusLane[3][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane19_strm1_data_valid    ( DownstreamStackBusLane[3][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane20_strm0_ready         ( DownstreamStackBusLane[3][20].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane20_strm0_cntl          ( DownstreamStackBusLane[3][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane20_strm0_data          ( DownstreamStackBusLane[3][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane20_strm0_data_valid    ( DownstreamStackBusLane[3][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane20_strm1_ready         ( DownstreamStackBusLane[3][20].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane20_strm1_cntl          ( DownstreamStackBusLane[3][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane20_strm1_data          ( DownstreamStackBusLane[3][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane20_strm1_data_valid    ( DownstreamStackBusLane[3][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane21_strm0_ready         ( DownstreamStackBusLane[3][21].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane21_strm0_cntl          ( DownstreamStackBusLane[3][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane21_strm0_data          ( DownstreamStackBusLane[3][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane21_strm0_data_valid    ( DownstreamStackBusLane[3][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane21_strm1_ready         ( DownstreamStackBusLane[3][21].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane21_strm1_cntl          ( DownstreamStackBusLane[3][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane21_strm1_data          ( DownstreamStackBusLane[3][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane21_strm1_data_valid    ( DownstreamStackBusLane[3][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane22_strm0_ready         ( DownstreamStackBusLane[3][22].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane22_strm0_cntl          ( DownstreamStackBusLane[3][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane22_strm0_data          ( DownstreamStackBusLane[3][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane22_strm0_data_valid    ( DownstreamStackBusLane[3][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane22_strm1_ready         ( DownstreamStackBusLane[3][22].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane22_strm1_cntl          ( DownstreamStackBusLane[3][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane22_strm1_data          ( DownstreamStackBusLane[3][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane22_strm1_data_valid    ( DownstreamStackBusLane[3][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane23_strm0_ready         ( DownstreamStackBusLane[3][23].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane23_strm0_cntl          ( DownstreamStackBusLane[3][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane23_strm0_data          ( DownstreamStackBusLane[3][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane23_strm0_data_valid    ( DownstreamStackBusLane[3][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane23_strm1_ready         ( DownstreamStackBusLane[3][23].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane23_strm1_cntl          ( DownstreamStackBusLane[3][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane23_strm1_data          ( DownstreamStackBusLane[3][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane23_strm1_data_valid    ( DownstreamStackBusLane[3][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane24_strm0_ready         ( DownstreamStackBusLane[3][24].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane24_strm0_cntl          ( DownstreamStackBusLane[3][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane24_strm0_data          ( DownstreamStackBusLane[3][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane24_strm0_data_valid    ( DownstreamStackBusLane[3][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane24_strm1_ready         ( DownstreamStackBusLane[3][24].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane24_strm1_cntl          ( DownstreamStackBusLane[3][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane24_strm1_data          ( DownstreamStackBusLane[3][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane24_strm1_data_valid    ( DownstreamStackBusLane[3][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane25_strm0_ready         ( DownstreamStackBusLane[3][25].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane25_strm0_cntl          ( DownstreamStackBusLane[3][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane25_strm0_data          ( DownstreamStackBusLane[3][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane25_strm0_data_valid    ( DownstreamStackBusLane[3][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane25_strm1_ready         ( DownstreamStackBusLane[3][25].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane25_strm1_cntl          ( DownstreamStackBusLane[3][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane25_strm1_data          ( DownstreamStackBusLane[3][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane25_strm1_data_valid    ( DownstreamStackBusLane[3][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane26_strm0_ready         ( DownstreamStackBusLane[3][26].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane26_strm0_cntl          ( DownstreamStackBusLane[3][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane26_strm0_data          ( DownstreamStackBusLane[3][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane26_strm0_data_valid    ( DownstreamStackBusLane[3][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane26_strm1_ready         ( DownstreamStackBusLane[3][26].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane26_strm1_cntl          ( DownstreamStackBusLane[3][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane26_strm1_data          ( DownstreamStackBusLane[3][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane26_strm1_data_valid    ( DownstreamStackBusLane[3][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane27_strm0_ready         ( DownstreamStackBusLane[3][27].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane27_strm0_cntl          ( DownstreamStackBusLane[3][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane27_strm0_data          ( DownstreamStackBusLane[3][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane27_strm0_data_valid    ( DownstreamStackBusLane[3][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane27_strm1_ready         ( DownstreamStackBusLane[3][27].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane27_strm1_cntl          ( DownstreamStackBusLane[3][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane27_strm1_data          ( DownstreamStackBusLane[3][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane27_strm1_data_valid    ( DownstreamStackBusLane[3][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane28_strm0_ready         ( DownstreamStackBusLane[3][28].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane28_strm0_cntl          ( DownstreamStackBusLane[3][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane28_strm0_data          ( DownstreamStackBusLane[3][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane28_strm0_data_valid    ( DownstreamStackBusLane[3][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane28_strm1_ready         ( DownstreamStackBusLane[3][28].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane28_strm1_cntl          ( DownstreamStackBusLane[3][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane28_strm1_data          ( DownstreamStackBusLane[3][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane28_strm1_data_valid    ( DownstreamStackBusLane[3][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane29_strm0_ready         ( DownstreamStackBusLane[3][29].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane29_strm0_cntl          ( DownstreamStackBusLane[3][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane29_strm0_data          ( DownstreamStackBusLane[3][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane29_strm0_data_valid    ( DownstreamStackBusLane[3][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane29_strm1_ready         ( DownstreamStackBusLane[3][29].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane29_strm1_cntl          ( DownstreamStackBusLane[3][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane29_strm1_data          ( DownstreamStackBusLane[3][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane29_strm1_data_valid    ( DownstreamStackBusLane[3][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane30_strm0_ready         ( DownstreamStackBusLane[3][30].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane30_strm0_cntl          ( DownstreamStackBusLane[3][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane30_strm0_data          ( DownstreamStackBusLane[3][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane30_strm0_data_valid    ( DownstreamStackBusLane[3][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane30_strm1_ready         ( DownstreamStackBusLane[3][30].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane30_strm1_cntl          ( DownstreamStackBusLane[3][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane30_strm1_data          ( DownstreamStackBusLane[3][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane30_strm1_data_valid    ( DownstreamStackBusLane[3][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane31_strm0_ready         ( DownstreamStackBusLane[3][31].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane31_strm0_cntl          ( DownstreamStackBusLane[3][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane31_strm0_data          ( DownstreamStackBusLane[3][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane31_strm0_data_valid    ( DownstreamStackBusLane[3][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane31_strm1_ready         ( DownstreamStackBusLane[3][31].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane31_strm1_cntl          ( DownstreamStackBusLane[3][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane31_strm1_data          ( DownstreamStackBusLane[3][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane31_strm1_data_valid    ( DownstreamStackBusLane[3][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane0_strm0_ready         ( DownstreamStackBusLane[4][0].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane0_strm0_cntl          ( DownstreamStackBusLane[4][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane0_strm0_data          ( DownstreamStackBusLane[4][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane0_strm0_data_valid    ( DownstreamStackBusLane[4][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane0_strm1_ready         ( DownstreamStackBusLane[4][0].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane0_strm1_cntl          ( DownstreamStackBusLane[4][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane0_strm1_data          ( DownstreamStackBusLane[4][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane0_strm1_data_valid    ( DownstreamStackBusLane[4][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane1_strm0_ready         ( DownstreamStackBusLane[4][1].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane1_strm0_cntl          ( DownstreamStackBusLane[4][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane1_strm0_data          ( DownstreamStackBusLane[4][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane1_strm0_data_valid    ( DownstreamStackBusLane[4][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane1_strm1_ready         ( DownstreamStackBusLane[4][1].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane1_strm1_cntl          ( DownstreamStackBusLane[4][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane1_strm1_data          ( DownstreamStackBusLane[4][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane1_strm1_data_valid    ( DownstreamStackBusLane[4][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane2_strm0_ready         ( DownstreamStackBusLane[4][2].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane2_strm0_cntl          ( DownstreamStackBusLane[4][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane2_strm0_data          ( DownstreamStackBusLane[4][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane2_strm0_data_valid    ( DownstreamStackBusLane[4][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane2_strm1_ready         ( DownstreamStackBusLane[4][2].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane2_strm1_cntl          ( DownstreamStackBusLane[4][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane2_strm1_data          ( DownstreamStackBusLane[4][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane2_strm1_data_valid    ( DownstreamStackBusLane[4][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane3_strm0_ready         ( DownstreamStackBusLane[4][3].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane3_strm0_cntl          ( DownstreamStackBusLane[4][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane3_strm0_data          ( DownstreamStackBusLane[4][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane3_strm0_data_valid    ( DownstreamStackBusLane[4][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane3_strm1_ready         ( DownstreamStackBusLane[4][3].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane3_strm1_cntl          ( DownstreamStackBusLane[4][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane3_strm1_data          ( DownstreamStackBusLane[4][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane3_strm1_data_valid    ( DownstreamStackBusLane[4][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane4_strm0_ready         ( DownstreamStackBusLane[4][4].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane4_strm0_cntl          ( DownstreamStackBusLane[4][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane4_strm0_data          ( DownstreamStackBusLane[4][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane4_strm0_data_valid    ( DownstreamStackBusLane[4][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane4_strm1_ready         ( DownstreamStackBusLane[4][4].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane4_strm1_cntl          ( DownstreamStackBusLane[4][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane4_strm1_data          ( DownstreamStackBusLane[4][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane4_strm1_data_valid    ( DownstreamStackBusLane[4][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane5_strm0_ready         ( DownstreamStackBusLane[4][5].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane5_strm0_cntl          ( DownstreamStackBusLane[4][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane5_strm0_data          ( DownstreamStackBusLane[4][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane5_strm0_data_valid    ( DownstreamStackBusLane[4][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane5_strm1_ready         ( DownstreamStackBusLane[4][5].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane5_strm1_cntl          ( DownstreamStackBusLane[4][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane5_strm1_data          ( DownstreamStackBusLane[4][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane5_strm1_data_valid    ( DownstreamStackBusLane[4][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane6_strm0_ready         ( DownstreamStackBusLane[4][6].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane6_strm0_cntl          ( DownstreamStackBusLane[4][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane6_strm0_data          ( DownstreamStackBusLane[4][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane6_strm0_data_valid    ( DownstreamStackBusLane[4][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane6_strm1_ready         ( DownstreamStackBusLane[4][6].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane6_strm1_cntl          ( DownstreamStackBusLane[4][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane6_strm1_data          ( DownstreamStackBusLane[4][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane6_strm1_data_valid    ( DownstreamStackBusLane[4][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane7_strm0_ready         ( DownstreamStackBusLane[4][7].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane7_strm0_cntl          ( DownstreamStackBusLane[4][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane7_strm0_data          ( DownstreamStackBusLane[4][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane7_strm0_data_valid    ( DownstreamStackBusLane[4][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane7_strm1_ready         ( DownstreamStackBusLane[4][7].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane7_strm1_cntl          ( DownstreamStackBusLane[4][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane7_strm1_data          ( DownstreamStackBusLane[4][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane7_strm1_data_valid    ( DownstreamStackBusLane[4][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane8_strm0_ready         ( DownstreamStackBusLane[4][8].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane8_strm0_cntl          ( DownstreamStackBusLane[4][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane8_strm0_data          ( DownstreamStackBusLane[4][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane8_strm0_data_valid    ( DownstreamStackBusLane[4][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane8_strm1_ready         ( DownstreamStackBusLane[4][8].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane8_strm1_cntl          ( DownstreamStackBusLane[4][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane8_strm1_data          ( DownstreamStackBusLane[4][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane8_strm1_data_valid    ( DownstreamStackBusLane[4][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane9_strm0_ready         ( DownstreamStackBusLane[4][9].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane9_strm0_cntl          ( DownstreamStackBusLane[4][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane9_strm0_data          ( DownstreamStackBusLane[4][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane9_strm0_data_valid    ( DownstreamStackBusLane[4][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane9_strm1_ready         ( DownstreamStackBusLane[4][9].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane9_strm1_cntl          ( DownstreamStackBusLane[4][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane9_strm1_data          ( DownstreamStackBusLane[4][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane9_strm1_data_valid    ( DownstreamStackBusLane[4][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane10_strm0_ready         ( DownstreamStackBusLane[4][10].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane10_strm0_cntl          ( DownstreamStackBusLane[4][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane10_strm0_data          ( DownstreamStackBusLane[4][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane10_strm0_data_valid    ( DownstreamStackBusLane[4][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane10_strm1_ready         ( DownstreamStackBusLane[4][10].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane10_strm1_cntl          ( DownstreamStackBusLane[4][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane10_strm1_data          ( DownstreamStackBusLane[4][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane10_strm1_data_valid    ( DownstreamStackBusLane[4][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane11_strm0_ready         ( DownstreamStackBusLane[4][11].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane11_strm0_cntl          ( DownstreamStackBusLane[4][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane11_strm0_data          ( DownstreamStackBusLane[4][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane11_strm0_data_valid    ( DownstreamStackBusLane[4][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane11_strm1_ready         ( DownstreamStackBusLane[4][11].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane11_strm1_cntl          ( DownstreamStackBusLane[4][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane11_strm1_data          ( DownstreamStackBusLane[4][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane11_strm1_data_valid    ( DownstreamStackBusLane[4][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane12_strm0_ready         ( DownstreamStackBusLane[4][12].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane12_strm0_cntl          ( DownstreamStackBusLane[4][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane12_strm0_data          ( DownstreamStackBusLane[4][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane12_strm0_data_valid    ( DownstreamStackBusLane[4][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane12_strm1_ready         ( DownstreamStackBusLane[4][12].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane12_strm1_cntl          ( DownstreamStackBusLane[4][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane12_strm1_data          ( DownstreamStackBusLane[4][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane12_strm1_data_valid    ( DownstreamStackBusLane[4][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane13_strm0_ready         ( DownstreamStackBusLane[4][13].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane13_strm0_cntl          ( DownstreamStackBusLane[4][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane13_strm0_data          ( DownstreamStackBusLane[4][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane13_strm0_data_valid    ( DownstreamStackBusLane[4][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane13_strm1_ready         ( DownstreamStackBusLane[4][13].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane13_strm1_cntl          ( DownstreamStackBusLane[4][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane13_strm1_data          ( DownstreamStackBusLane[4][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane13_strm1_data_valid    ( DownstreamStackBusLane[4][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane14_strm0_ready         ( DownstreamStackBusLane[4][14].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane14_strm0_cntl          ( DownstreamStackBusLane[4][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane14_strm0_data          ( DownstreamStackBusLane[4][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane14_strm0_data_valid    ( DownstreamStackBusLane[4][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane14_strm1_ready         ( DownstreamStackBusLane[4][14].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane14_strm1_cntl          ( DownstreamStackBusLane[4][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane14_strm1_data          ( DownstreamStackBusLane[4][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane14_strm1_data_valid    ( DownstreamStackBusLane[4][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane15_strm0_ready         ( DownstreamStackBusLane[4][15].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane15_strm0_cntl          ( DownstreamStackBusLane[4][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane15_strm0_data          ( DownstreamStackBusLane[4][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane15_strm0_data_valid    ( DownstreamStackBusLane[4][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane15_strm1_ready         ( DownstreamStackBusLane[4][15].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane15_strm1_cntl          ( DownstreamStackBusLane[4][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane15_strm1_data          ( DownstreamStackBusLane[4][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane15_strm1_data_valid    ( DownstreamStackBusLane[4][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane16_strm0_ready         ( DownstreamStackBusLane[4][16].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane16_strm0_cntl          ( DownstreamStackBusLane[4][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane16_strm0_data          ( DownstreamStackBusLane[4][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane16_strm0_data_valid    ( DownstreamStackBusLane[4][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane16_strm1_ready         ( DownstreamStackBusLane[4][16].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane16_strm1_cntl          ( DownstreamStackBusLane[4][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane16_strm1_data          ( DownstreamStackBusLane[4][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane16_strm1_data_valid    ( DownstreamStackBusLane[4][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane17_strm0_ready         ( DownstreamStackBusLane[4][17].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane17_strm0_cntl          ( DownstreamStackBusLane[4][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane17_strm0_data          ( DownstreamStackBusLane[4][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane17_strm0_data_valid    ( DownstreamStackBusLane[4][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane17_strm1_ready         ( DownstreamStackBusLane[4][17].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane17_strm1_cntl          ( DownstreamStackBusLane[4][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane17_strm1_data          ( DownstreamStackBusLane[4][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane17_strm1_data_valid    ( DownstreamStackBusLane[4][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane18_strm0_ready         ( DownstreamStackBusLane[4][18].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane18_strm0_cntl          ( DownstreamStackBusLane[4][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane18_strm0_data          ( DownstreamStackBusLane[4][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane18_strm0_data_valid    ( DownstreamStackBusLane[4][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane18_strm1_ready         ( DownstreamStackBusLane[4][18].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane18_strm1_cntl          ( DownstreamStackBusLane[4][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane18_strm1_data          ( DownstreamStackBusLane[4][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane18_strm1_data_valid    ( DownstreamStackBusLane[4][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane19_strm0_ready         ( DownstreamStackBusLane[4][19].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane19_strm0_cntl          ( DownstreamStackBusLane[4][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane19_strm0_data          ( DownstreamStackBusLane[4][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane19_strm0_data_valid    ( DownstreamStackBusLane[4][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane19_strm1_ready         ( DownstreamStackBusLane[4][19].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane19_strm1_cntl          ( DownstreamStackBusLane[4][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane19_strm1_data          ( DownstreamStackBusLane[4][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane19_strm1_data_valid    ( DownstreamStackBusLane[4][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane20_strm0_ready         ( DownstreamStackBusLane[4][20].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane20_strm0_cntl          ( DownstreamStackBusLane[4][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane20_strm0_data          ( DownstreamStackBusLane[4][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane20_strm0_data_valid    ( DownstreamStackBusLane[4][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane20_strm1_ready         ( DownstreamStackBusLane[4][20].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane20_strm1_cntl          ( DownstreamStackBusLane[4][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane20_strm1_data          ( DownstreamStackBusLane[4][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane20_strm1_data_valid    ( DownstreamStackBusLane[4][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane21_strm0_ready         ( DownstreamStackBusLane[4][21].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane21_strm0_cntl          ( DownstreamStackBusLane[4][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane21_strm0_data          ( DownstreamStackBusLane[4][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane21_strm0_data_valid    ( DownstreamStackBusLane[4][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane21_strm1_ready         ( DownstreamStackBusLane[4][21].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane21_strm1_cntl          ( DownstreamStackBusLane[4][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane21_strm1_data          ( DownstreamStackBusLane[4][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane21_strm1_data_valid    ( DownstreamStackBusLane[4][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane22_strm0_ready         ( DownstreamStackBusLane[4][22].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane22_strm0_cntl          ( DownstreamStackBusLane[4][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane22_strm0_data          ( DownstreamStackBusLane[4][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane22_strm0_data_valid    ( DownstreamStackBusLane[4][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane22_strm1_ready         ( DownstreamStackBusLane[4][22].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane22_strm1_cntl          ( DownstreamStackBusLane[4][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane22_strm1_data          ( DownstreamStackBusLane[4][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane22_strm1_data_valid    ( DownstreamStackBusLane[4][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane23_strm0_ready         ( DownstreamStackBusLane[4][23].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane23_strm0_cntl          ( DownstreamStackBusLane[4][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane23_strm0_data          ( DownstreamStackBusLane[4][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane23_strm0_data_valid    ( DownstreamStackBusLane[4][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane23_strm1_ready         ( DownstreamStackBusLane[4][23].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane23_strm1_cntl          ( DownstreamStackBusLane[4][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane23_strm1_data          ( DownstreamStackBusLane[4][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane23_strm1_data_valid    ( DownstreamStackBusLane[4][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane24_strm0_ready         ( DownstreamStackBusLane[4][24].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane24_strm0_cntl          ( DownstreamStackBusLane[4][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane24_strm0_data          ( DownstreamStackBusLane[4][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane24_strm0_data_valid    ( DownstreamStackBusLane[4][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane24_strm1_ready         ( DownstreamStackBusLane[4][24].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane24_strm1_cntl          ( DownstreamStackBusLane[4][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane24_strm1_data          ( DownstreamStackBusLane[4][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane24_strm1_data_valid    ( DownstreamStackBusLane[4][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane25_strm0_ready         ( DownstreamStackBusLane[4][25].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane25_strm0_cntl          ( DownstreamStackBusLane[4][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane25_strm0_data          ( DownstreamStackBusLane[4][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane25_strm0_data_valid    ( DownstreamStackBusLane[4][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane25_strm1_ready         ( DownstreamStackBusLane[4][25].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane25_strm1_cntl          ( DownstreamStackBusLane[4][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane25_strm1_data          ( DownstreamStackBusLane[4][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane25_strm1_data_valid    ( DownstreamStackBusLane[4][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane26_strm0_ready         ( DownstreamStackBusLane[4][26].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane26_strm0_cntl          ( DownstreamStackBusLane[4][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane26_strm0_data          ( DownstreamStackBusLane[4][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane26_strm0_data_valid    ( DownstreamStackBusLane[4][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane26_strm1_ready         ( DownstreamStackBusLane[4][26].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane26_strm1_cntl          ( DownstreamStackBusLane[4][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane26_strm1_data          ( DownstreamStackBusLane[4][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane26_strm1_data_valid    ( DownstreamStackBusLane[4][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane27_strm0_ready         ( DownstreamStackBusLane[4][27].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane27_strm0_cntl          ( DownstreamStackBusLane[4][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane27_strm0_data          ( DownstreamStackBusLane[4][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane27_strm0_data_valid    ( DownstreamStackBusLane[4][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane27_strm1_ready         ( DownstreamStackBusLane[4][27].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane27_strm1_cntl          ( DownstreamStackBusLane[4][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane27_strm1_data          ( DownstreamStackBusLane[4][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane27_strm1_data_valid    ( DownstreamStackBusLane[4][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane28_strm0_ready         ( DownstreamStackBusLane[4][28].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane28_strm0_cntl          ( DownstreamStackBusLane[4][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane28_strm0_data          ( DownstreamStackBusLane[4][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane28_strm0_data_valid    ( DownstreamStackBusLane[4][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane28_strm1_ready         ( DownstreamStackBusLane[4][28].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane28_strm1_cntl          ( DownstreamStackBusLane[4][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane28_strm1_data          ( DownstreamStackBusLane[4][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane28_strm1_data_valid    ( DownstreamStackBusLane[4][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane29_strm0_ready         ( DownstreamStackBusLane[4][29].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane29_strm0_cntl          ( DownstreamStackBusLane[4][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane29_strm0_data          ( DownstreamStackBusLane[4][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane29_strm0_data_valid    ( DownstreamStackBusLane[4][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane29_strm1_ready         ( DownstreamStackBusLane[4][29].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane29_strm1_cntl          ( DownstreamStackBusLane[4][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane29_strm1_data          ( DownstreamStackBusLane[4][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane29_strm1_data_valid    ( DownstreamStackBusLane[4][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane30_strm0_ready         ( DownstreamStackBusLane[4][30].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane30_strm0_cntl          ( DownstreamStackBusLane[4][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane30_strm0_data          ( DownstreamStackBusLane[4][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane30_strm0_data_valid    ( DownstreamStackBusLane[4][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane30_strm1_ready         ( DownstreamStackBusLane[4][30].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane30_strm1_cntl          ( DownstreamStackBusLane[4][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane30_strm1_data          ( DownstreamStackBusLane[4][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane30_strm1_data_valid    ( DownstreamStackBusLane[4][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 4, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane31_strm0_ready         ( DownstreamStackBusLane[4][31].pe__std__lane_strm0_ready              ),      
        .std__pe4__lane31_strm0_cntl          ( DownstreamStackBusLane[4][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe4__lane31_strm0_data          ( DownstreamStackBusLane[4][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe4__lane31_strm0_data_valid    ( DownstreamStackBusLane[4][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__std__lane31_strm1_ready         ( DownstreamStackBusLane[4][31].pe__std__lane_strm1_ready              ),      
        .std__pe4__lane31_strm1_cntl          ( DownstreamStackBusLane[4][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe4__lane31_strm1_data          ( DownstreamStackBusLane[4][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe4__lane31_strm1_data_valid    ( DownstreamStackBusLane[4][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane0_strm0_ready         ( DownstreamStackBusLane[5][0].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane0_strm0_cntl          ( DownstreamStackBusLane[5][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane0_strm0_data          ( DownstreamStackBusLane[5][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane0_strm0_data_valid    ( DownstreamStackBusLane[5][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane0_strm1_ready         ( DownstreamStackBusLane[5][0].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane0_strm1_cntl          ( DownstreamStackBusLane[5][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane0_strm1_data          ( DownstreamStackBusLane[5][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane0_strm1_data_valid    ( DownstreamStackBusLane[5][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane1_strm0_ready         ( DownstreamStackBusLane[5][1].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane1_strm0_cntl          ( DownstreamStackBusLane[5][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane1_strm0_data          ( DownstreamStackBusLane[5][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane1_strm0_data_valid    ( DownstreamStackBusLane[5][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane1_strm1_ready         ( DownstreamStackBusLane[5][1].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane1_strm1_cntl          ( DownstreamStackBusLane[5][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane1_strm1_data          ( DownstreamStackBusLane[5][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane1_strm1_data_valid    ( DownstreamStackBusLane[5][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane2_strm0_ready         ( DownstreamStackBusLane[5][2].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane2_strm0_cntl          ( DownstreamStackBusLane[5][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane2_strm0_data          ( DownstreamStackBusLane[5][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane2_strm0_data_valid    ( DownstreamStackBusLane[5][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane2_strm1_ready         ( DownstreamStackBusLane[5][2].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane2_strm1_cntl          ( DownstreamStackBusLane[5][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane2_strm1_data          ( DownstreamStackBusLane[5][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane2_strm1_data_valid    ( DownstreamStackBusLane[5][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane3_strm0_ready         ( DownstreamStackBusLane[5][3].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane3_strm0_cntl          ( DownstreamStackBusLane[5][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane3_strm0_data          ( DownstreamStackBusLane[5][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane3_strm0_data_valid    ( DownstreamStackBusLane[5][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane3_strm1_ready         ( DownstreamStackBusLane[5][3].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane3_strm1_cntl          ( DownstreamStackBusLane[5][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane3_strm1_data          ( DownstreamStackBusLane[5][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane3_strm1_data_valid    ( DownstreamStackBusLane[5][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane4_strm0_ready         ( DownstreamStackBusLane[5][4].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane4_strm0_cntl          ( DownstreamStackBusLane[5][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane4_strm0_data          ( DownstreamStackBusLane[5][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane4_strm0_data_valid    ( DownstreamStackBusLane[5][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane4_strm1_ready         ( DownstreamStackBusLane[5][4].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane4_strm1_cntl          ( DownstreamStackBusLane[5][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane4_strm1_data          ( DownstreamStackBusLane[5][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane4_strm1_data_valid    ( DownstreamStackBusLane[5][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane5_strm0_ready         ( DownstreamStackBusLane[5][5].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane5_strm0_cntl          ( DownstreamStackBusLane[5][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane5_strm0_data          ( DownstreamStackBusLane[5][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane5_strm0_data_valid    ( DownstreamStackBusLane[5][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane5_strm1_ready         ( DownstreamStackBusLane[5][5].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane5_strm1_cntl          ( DownstreamStackBusLane[5][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane5_strm1_data          ( DownstreamStackBusLane[5][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane5_strm1_data_valid    ( DownstreamStackBusLane[5][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane6_strm0_ready         ( DownstreamStackBusLane[5][6].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane6_strm0_cntl          ( DownstreamStackBusLane[5][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane6_strm0_data          ( DownstreamStackBusLane[5][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane6_strm0_data_valid    ( DownstreamStackBusLane[5][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane6_strm1_ready         ( DownstreamStackBusLane[5][6].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane6_strm1_cntl          ( DownstreamStackBusLane[5][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane6_strm1_data          ( DownstreamStackBusLane[5][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane6_strm1_data_valid    ( DownstreamStackBusLane[5][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane7_strm0_ready         ( DownstreamStackBusLane[5][7].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane7_strm0_cntl          ( DownstreamStackBusLane[5][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane7_strm0_data          ( DownstreamStackBusLane[5][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane7_strm0_data_valid    ( DownstreamStackBusLane[5][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane7_strm1_ready         ( DownstreamStackBusLane[5][7].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane7_strm1_cntl          ( DownstreamStackBusLane[5][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane7_strm1_data          ( DownstreamStackBusLane[5][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane7_strm1_data_valid    ( DownstreamStackBusLane[5][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane8_strm0_ready         ( DownstreamStackBusLane[5][8].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane8_strm0_cntl          ( DownstreamStackBusLane[5][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane8_strm0_data          ( DownstreamStackBusLane[5][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane8_strm0_data_valid    ( DownstreamStackBusLane[5][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane8_strm1_ready         ( DownstreamStackBusLane[5][8].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane8_strm1_cntl          ( DownstreamStackBusLane[5][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane8_strm1_data          ( DownstreamStackBusLane[5][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane8_strm1_data_valid    ( DownstreamStackBusLane[5][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane9_strm0_ready         ( DownstreamStackBusLane[5][9].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane9_strm0_cntl          ( DownstreamStackBusLane[5][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane9_strm0_data          ( DownstreamStackBusLane[5][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane9_strm0_data_valid    ( DownstreamStackBusLane[5][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane9_strm1_ready         ( DownstreamStackBusLane[5][9].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane9_strm1_cntl          ( DownstreamStackBusLane[5][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane9_strm1_data          ( DownstreamStackBusLane[5][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane9_strm1_data_valid    ( DownstreamStackBusLane[5][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane10_strm0_ready         ( DownstreamStackBusLane[5][10].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane10_strm0_cntl          ( DownstreamStackBusLane[5][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane10_strm0_data          ( DownstreamStackBusLane[5][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane10_strm0_data_valid    ( DownstreamStackBusLane[5][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane10_strm1_ready         ( DownstreamStackBusLane[5][10].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane10_strm1_cntl          ( DownstreamStackBusLane[5][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane10_strm1_data          ( DownstreamStackBusLane[5][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane10_strm1_data_valid    ( DownstreamStackBusLane[5][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane11_strm0_ready         ( DownstreamStackBusLane[5][11].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane11_strm0_cntl          ( DownstreamStackBusLane[5][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane11_strm0_data          ( DownstreamStackBusLane[5][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane11_strm0_data_valid    ( DownstreamStackBusLane[5][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane11_strm1_ready         ( DownstreamStackBusLane[5][11].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane11_strm1_cntl          ( DownstreamStackBusLane[5][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane11_strm1_data          ( DownstreamStackBusLane[5][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane11_strm1_data_valid    ( DownstreamStackBusLane[5][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane12_strm0_ready         ( DownstreamStackBusLane[5][12].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane12_strm0_cntl          ( DownstreamStackBusLane[5][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane12_strm0_data          ( DownstreamStackBusLane[5][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane12_strm0_data_valid    ( DownstreamStackBusLane[5][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane12_strm1_ready         ( DownstreamStackBusLane[5][12].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane12_strm1_cntl          ( DownstreamStackBusLane[5][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane12_strm1_data          ( DownstreamStackBusLane[5][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane12_strm1_data_valid    ( DownstreamStackBusLane[5][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane13_strm0_ready         ( DownstreamStackBusLane[5][13].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane13_strm0_cntl          ( DownstreamStackBusLane[5][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane13_strm0_data          ( DownstreamStackBusLane[5][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane13_strm0_data_valid    ( DownstreamStackBusLane[5][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane13_strm1_ready         ( DownstreamStackBusLane[5][13].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane13_strm1_cntl          ( DownstreamStackBusLane[5][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane13_strm1_data          ( DownstreamStackBusLane[5][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane13_strm1_data_valid    ( DownstreamStackBusLane[5][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane14_strm0_ready         ( DownstreamStackBusLane[5][14].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane14_strm0_cntl          ( DownstreamStackBusLane[5][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane14_strm0_data          ( DownstreamStackBusLane[5][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane14_strm0_data_valid    ( DownstreamStackBusLane[5][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane14_strm1_ready         ( DownstreamStackBusLane[5][14].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane14_strm1_cntl          ( DownstreamStackBusLane[5][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane14_strm1_data          ( DownstreamStackBusLane[5][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane14_strm1_data_valid    ( DownstreamStackBusLane[5][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane15_strm0_ready         ( DownstreamStackBusLane[5][15].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane15_strm0_cntl          ( DownstreamStackBusLane[5][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane15_strm0_data          ( DownstreamStackBusLane[5][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane15_strm0_data_valid    ( DownstreamStackBusLane[5][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane15_strm1_ready         ( DownstreamStackBusLane[5][15].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane15_strm1_cntl          ( DownstreamStackBusLane[5][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane15_strm1_data          ( DownstreamStackBusLane[5][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane15_strm1_data_valid    ( DownstreamStackBusLane[5][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane16_strm0_ready         ( DownstreamStackBusLane[5][16].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane16_strm0_cntl          ( DownstreamStackBusLane[5][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane16_strm0_data          ( DownstreamStackBusLane[5][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane16_strm0_data_valid    ( DownstreamStackBusLane[5][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane16_strm1_ready         ( DownstreamStackBusLane[5][16].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane16_strm1_cntl          ( DownstreamStackBusLane[5][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane16_strm1_data          ( DownstreamStackBusLane[5][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane16_strm1_data_valid    ( DownstreamStackBusLane[5][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane17_strm0_ready         ( DownstreamStackBusLane[5][17].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane17_strm0_cntl          ( DownstreamStackBusLane[5][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane17_strm0_data          ( DownstreamStackBusLane[5][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane17_strm0_data_valid    ( DownstreamStackBusLane[5][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane17_strm1_ready         ( DownstreamStackBusLane[5][17].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane17_strm1_cntl          ( DownstreamStackBusLane[5][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane17_strm1_data          ( DownstreamStackBusLane[5][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane17_strm1_data_valid    ( DownstreamStackBusLane[5][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane18_strm0_ready         ( DownstreamStackBusLane[5][18].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane18_strm0_cntl          ( DownstreamStackBusLane[5][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane18_strm0_data          ( DownstreamStackBusLane[5][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane18_strm0_data_valid    ( DownstreamStackBusLane[5][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane18_strm1_ready         ( DownstreamStackBusLane[5][18].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane18_strm1_cntl          ( DownstreamStackBusLane[5][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane18_strm1_data          ( DownstreamStackBusLane[5][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane18_strm1_data_valid    ( DownstreamStackBusLane[5][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane19_strm0_ready         ( DownstreamStackBusLane[5][19].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane19_strm0_cntl          ( DownstreamStackBusLane[5][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane19_strm0_data          ( DownstreamStackBusLane[5][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane19_strm0_data_valid    ( DownstreamStackBusLane[5][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane19_strm1_ready         ( DownstreamStackBusLane[5][19].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane19_strm1_cntl          ( DownstreamStackBusLane[5][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane19_strm1_data          ( DownstreamStackBusLane[5][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane19_strm1_data_valid    ( DownstreamStackBusLane[5][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane20_strm0_ready         ( DownstreamStackBusLane[5][20].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane20_strm0_cntl          ( DownstreamStackBusLane[5][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane20_strm0_data          ( DownstreamStackBusLane[5][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane20_strm0_data_valid    ( DownstreamStackBusLane[5][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane20_strm1_ready         ( DownstreamStackBusLane[5][20].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane20_strm1_cntl          ( DownstreamStackBusLane[5][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane20_strm1_data          ( DownstreamStackBusLane[5][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane20_strm1_data_valid    ( DownstreamStackBusLane[5][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane21_strm0_ready         ( DownstreamStackBusLane[5][21].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane21_strm0_cntl          ( DownstreamStackBusLane[5][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane21_strm0_data          ( DownstreamStackBusLane[5][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane21_strm0_data_valid    ( DownstreamStackBusLane[5][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane21_strm1_ready         ( DownstreamStackBusLane[5][21].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane21_strm1_cntl          ( DownstreamStackBusLane[5][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane21_strm1_data          ( DownstreamStackBusLane[5][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane21_strm1_data_valid    ( DownstreamStackBusLane[5][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane22_strm0_ready         ( DownstreamStackBusLane[5][22].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane22_strm0_cntl          ( DownstreamStackBusLane[5][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane22_strm0_data          ( DownstreamStackBusLane[5][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane22_strm0_data_valid    ( DownstreamStackBusLane[5][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane22_strm1_ready         ( DownstreamStackBusLane[5][22].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane22_strm1_cntl          ( DownstreamStackBusLane[5][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane22_strm1_data          ( DownstreamStackBusLane[5][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane22_strm1_data_valid    ( DownstreamStackBusLane[5][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane23_strm0_ready         ( DownstreamStackBusLane[5][23].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane23_strm0_cntl          ( DownstreamStackBusLane[5][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane23_strm0_data          ( DownstreamStackBusLane[5][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane23_strm0_data_valid    ( DownstreamStackBusLane[5][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane23_strm1_ready         ( DownstreamStackBusLane[5][23].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane23_strm1_cntl          ( DownstreamStackBusLane[5][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane23_strm1_data          ( DownstreamStackBusLane[5][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane23_strm1_data_valid    ( DownstreamStackBusLane[5][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane24_strm0_ready         ( DownstreamStackBusLane[5][24].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane24_strm0_cntl          ( DownstreamStackBusLane[5][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane24_strm0_data          ( DownstreamStackBusLane[5][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane24_strm0_data_valid    ( DownstreamStackBusLane[5][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane24_strm1_ready         ( DownstreamStackBusLane[5][24].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane24_strm1_cntl          ( DownstreamStackBusLane[5][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane24_strm1_data          ( DownstreamStackBusLane[5][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane24_strm1_data_valid    ( DownstreamStackBusLane[5][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane25_strm0_ready         ( DownstreamStackBusLane[5][25].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane25_strm0_cntl          ( DownstreamStackBusLane[5][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane25_strm0_data          ( DownstreamStackBusLane[5][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane25_strm0_data_valid    ( DownstreamStackBusLane[5][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane25_strm1_ready         ( DownstreamStackBusLane[5][25].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane25_strm1_cntl          ( DownstreamStackBusLane[5][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane25_strm1_data          ( DownstreamStackBusLane[5][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane25_strm1_data_valid    ( DownstreamStackBusLane[5][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane26_strm0_ready         ( DownstreamStackBusLane[5][26].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane26_strm0_cntl          ( DownstreamStackBusLane[5][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane26_strm0_data          ( DownstreamStackBusLane[5][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane26_strm0_data_valid    ( DownstreamStackBusLane[5][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane26_strm1_ready         ( DownstreamStackBusLane[5][26].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane26_strm1_cntl          ( DownstreamStackBusLane[5][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane26_strm1_data          ( DownstreamStackBusLane[5][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane26_strm1_data_valid    ( DownstreamStackBusLane[5][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane27_strm0_ready         ( DownstreamStackBusLane[5][27].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane27_strm0_cntl          ( DownstreamStackBusLane[5][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane27_strm0_data          ( DownstreamStackBusLane[5][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane27_strm0_data_valid    ( DownstreamStackBusLane[5][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane27_strm1_ready         ( DownstreamStackBusLane[5][27].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane27_strm1_cntl          ( DownstreamStackBusLane[5][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane27_strm1_data          ( DownstreamStackBusLane[5][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane27_strm1_data_valid    ( DownstreamStackBusLane[5][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane28_strm0_ready         ( DownstreamStackBusLane[5][28].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane28_strm0_cntl          ( DownstreamStackBusLane[5][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane28_strm0_data          ( DownstreamStackBusLane[5][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane28_strm0_data_valid    ( DownstreamStackBusLane[5][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane28_strm1_ready         ( DownstreamStackBusLane[5][28].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane28_strm1_cntl          ( DownstreamStackBusLane[5][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane28_strm1_data          ( DownstreamStackBusLane[5][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane28_strm1_data_valid    ( DownstreamStackBusLane[5][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane29_strm0_ready         ( DownstreamStackBusLane[5][29].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane29_strm0_cntl          ( DownstreamStackBusLane[5][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane29_strm0_data          ( DownstreamStackBusLane[5][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane29_strm0_data_valid    ( DownstreamStackBusLane[5][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane29_strm1_ready         ( DownstreamStackBusLane[5][29].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane29_strm1_cntl          ( DownstreamStackBusLane[5][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane29_strm1_data          ( DownstreamStackBusLane[5][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane29_strm1_data_valid    ( DownstreamStackBusLane[5][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane30_strm0_ready         ( DownstreamStackBusLane[5][30].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane30_strm0_cntl          ( DownstreamStackBusLane[5][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane30_strm0_data          ( DownstreamStackBusLane[5][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane30_strm0_data_valid    ( DownstreamStackBusLane[5][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane30_strm1_ready         ( DownstreamStackBusLane[5][30].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane30_strm1_cntl          ( DownstreamStackBusLane[5][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane30_strm1_data          ( DownstreamStackBusLane[5][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane30_strm1_data_valid    ( DownstreamStackBusLane[5][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 5, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane31_strm0_ready         ( DownstreamStackBusLane[5][31].pe__std__lane_strm0_ready              ),      
        .std__pe5__lane31_strm0_cntl          ( DownstreamStackBusLane[5][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe5__lane31_strm0_data          ( DownstreamStackBusLane[5][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe5__lane31_strm0_data_valid    ( DownstreamStackBusLane[5][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__std__lane31_strm1_ready         ( DownstreamStackBusLane[5][31].pe__std__lane_strm1_ready              ),      
        .std__pe5__lane31_strm1_cntl          ( DownstreamStackBusLane[5][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe5__lane31_strm1_data          ( DownstreamStackBusLane[5][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe5__lane31_strm1_data_valid    ( DownstreamStackBusLane[5][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane0_strm0_ready         ( DownstreamStackBusLane[6][0].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane0_strm0_cntl          ( DownstreamStackBusLane[6][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane0_strm0_data          ( DownstreamStackBusLane[6][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane0_strm0_data_valid    ( DownstreamStackBusLane[6][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane0_strm1_ready         ( DownstreamStackBusLane[6][0].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane0_strm1_cntl          ( DownstreamStackBusLane[6][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane0_strm1_data          ( DownstreamStackBusLane[6][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane0_strm1_data_valid    ( DownstreamStackBusLane[6][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane1_strm0_ready         ( DownstreamStackBusLane[6][1].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane1_strm0_cntl          ( DownstreamStackBusLane[6][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane1_strm0_data          ( DownstreamStackBusLane[6][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane1_strm0_data_valid    ( DownstreamStackBusLane[6][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane1_strm1_ready         ( DownstreamStackBusLane[6][1].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane1_strm1_cntl          ( DownstreamStackBusLane[6][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane1_strm1_data          ( DownstreamStackBusLane[6][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane1_strm1_data_valid    ( DownstreamStackBusLane[6][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane2_strm0_ready         ( DownstreamStackBusLane[6][2].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane2_strm0_cntl          ( DownstreamStackBusLane[6][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane2_strm0_data          ( DownstreamStackBusLane[6][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane2_strm0_data_valid    ( DownstreamStackBusLane[6][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane2_strm1_ready         ( DownstreamStackBusLane[6][2].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane2_strm1_cntl          ( DownstreamStackBusLane[6][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane2_strm1_data          ( DownstreamStackBusLane[6][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane2_strm1_data_valid    ( DownstreamStackBusLane[6][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane3_strm0_ready         ( DownstreamStackBusLane[6][3].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane3_strm0_cntl          ( DownstreamStackBusLane[6][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane3_strm0_data          ( DownstreamStackBusLane[6][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane3_strm0_data_valid    ( DownstreamStackBusLane[6][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane3_strm1_ready         ( DownstreamStackBusLane[6][3].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane3_strm1_cntl          ( DownstreamStackBusLane[6][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane3_strm1_data          ( DownstreamStackBusLane[6][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane3_strm1_data_valid    ( DownstreamStackBusLane[6][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane4_strm0_ready         ( DownstreamStackBusLane[6][4].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane4_strm0_cntl          ( DownstreamStackBusLane[6][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane4_strm0_data          ( DownstreamStackBusLane[6][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane4_strm0_data_valid    ( DownstreamStackBusLane[6][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane4_strm1_ready         ( DownstreamStackBusLane[6][4].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane4_strm1_cntl          ( DownstreamStackBusLane[6][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane4_strm1_data          ( DownstreamStackBusLane[6][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane4_strm1_data_valid    ( DownstreamStackBusLane[6][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane5_strm0_ready         ( DownstreamStackBusLane[6][5].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane5_strm0_cntl          ( DownstreamStackBusLane[6][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane5_strm0_data          ( DownstreamStackBusLane[6][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane5_strm0_data_valid    ( DownstreamStackBusLane[6][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane5_strm1_ready         ( DownstreamStackBusLane[6][5].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane5_strm1_cntl          ( DownstreamStackBusLane[6][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane5_strm1_data          ( DownstreamStackBusLane[6][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane5_strm1_data_valid    ( DownstreamStackBusLane[6][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane6_strm0_ready         ( DownstreamStackBusLane[6][6].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane6_strm0_cntl          ( DownstreamStackBusLane[6][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane6_strm0_data          ( DownstreamStackBusLane[6][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane6_strm0_data_valid    ( DownstreamStackBusLane[6][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane6_strm1_ready         ( DownstreamStackBusLane[6][6].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane6_strm1_cntl          ( DownstreamStackBusLane[6][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane6_strm1_data          ( DownstreamStackBusLane[6][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane6_strm1_data_valid    ( DownstreamStackBusLane[6][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane7_strm0_ready         ( DownstreamStackBusLane[6][7].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane7_strm0_cntl          ( DownstreamStackBusLane[6][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane7_strm0_data          ( DownstreamStackBusLane[6][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane7_strm0_data_valid    ( DownstreamStackBusLane[6][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane7_strm1_ready         ( DownstreamStackBusLane[6][7].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane7_strm1_cntl          ( DownstreamStackBusLane[6][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane7_strm1_data          ( DownstreamStackBusLane[6][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane7_strm1_data_valid    ( DownstreamStackBusLane[6][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane8_strm0_ready         ( DownstreamStackBusLane[6][8].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane8_strm0_cntl          ( DownstreamStackBusLane[6][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane8_strm0_data          ( DownstreamStackBusLane[6][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane8_strm0_data_valid    ( DownstreamStackBusLane[6][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane8_strm1_ready         ( DownstreamStackBusLane[6][8].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane8_strm1_cntl          ( DownstreamStackBusLane[6][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane8_strm1_data          ( DownstreamStackBusLane[6][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane8_strm1_data_valid    ( DownstreamStackBusLane[6][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane9_strm0_ready         ( DownstreamStackBusLane[6][9].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane9_strm0_cntl          ( DownstreamStackBusLane[6][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane9_strm0_data          ( DownstreamStackBusLane[6][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane9_strm0_data_valid    ( DownstreamStackBusLane[6][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane9_strm1_ready         ( DownstreamStackBusLane[6][9].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane9_strm1_cntl          ( DownstreamStackBusLane[6][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane9_strm1_data          ( DownstreamStackBusLane[6][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane9_strm1_data_valid    ( DownstreamStackBusLane[6][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane10_strm0_ready         ( DownstreamStackBusLane[6][10].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane10_strm0_cntl          ( DownstreamStackBusLane[6][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane10_strm0_data          ( DownstreamStackBusLane[6][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane10_strm0_data_valid    ( DownstreamStackBusLane[6][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane10_strm1_ready         ( DownstreamStackBusLane[6][10].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane10_strm1_cntl          ( DownstreamStackBusLane[6][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane10_strm1_data          ( DownstreamStackBusLane[6][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane10_strm1_data_valid    ( DownstreamStackBusLane[6][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane11_strm0_ready         ( DownstreamStackBusLane[6][11].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane11_strm0_cntl          ( DownstreamStackBusLane[6][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane11_strm0_data          ( DownstreamStackBusLane[6][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane11_strm0_data_valid    ( DownstreamStackBusLane[6][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane11_strm1_ready         ( DownstreamStackBusLane[6][11].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane11_strm1_cntl          ( DownstreamStackBusLane[6][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane11_strm1_data          ( DownstreamStackBusLane[6][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane11_strm1_data_valid    ( DownstreamStackBusLane[6][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane12_strm0_ready         ( DownstreamStackBusLane[6][12].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane12_strm0_cntl          ( DownstreamStackBusLane[6][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane12_strm0_data          ( DownstreamStackBusLane[6][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane12_strm0_data_valid    ( DownstreamStackBusLane[6][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane12_strm1_ready         ( DownstreamStackBusLane[6][12].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane12_strm1_cntl          ( DownstreamStackBusLane[6][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane12_strm1_data          ( DownstreamStackBusLane[6][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane12_strm1_data_valid    ( DownstreamStackBusLane[6][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane13_strm0_ready         ( DownstreamStackBusLane[6][13].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane13_strm0_cntl          ( DownstreamStackBusLane[6][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane13_strm0_data          ( DownstreamStackBusLane[6][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane13_strm0_data_valid    ( DownstreamStackBusLane[6][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane13_strm1_ready         ( DownstreamStackBusLane[6][13].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane13_strm1_cntl          ( DownstreamStackBusLane[6][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane13_strm1_data          ( DownstreamStackBusLane[6][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane13_strm1_data_valid    ( DownstreamStackBusLane[6][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane14_strm0_ready         ( DownstreamStackBusLane[6][14].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane14_strm0_cntl          ( DownstreamStackBusLane[6][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane14_strm0_data          ( DownstreamStackBusLane[6][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane14_strm0_data_valid    ( DownstreamStackBusLane[6][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane14_strm1_ready         ( DownstreamStackBusLane[6][14].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane14_strm1_cntl          ( DownstreamStackBusLane[6][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane14_strm1_data          ( DownstreamStackBusLane[6][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane14_strm1_data_valid    ( DownstreamStackBusLane[6][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane15_strm0_ready         ( DownstreamStackBusLane[6][15].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane15_strm0_cntl          ( DownstreamStackBusLane[6][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane15_strm0_data          ( DownstreamStackBusLane[6][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane15_strm0_data_valid    ( DownstreamStackBusLane[6][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane15_strm1_ready         ( DownstreamStackBusLane[6][15].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane15_strm1_cntl          ( DownstreamStackBusLane[6][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane15_strm1_data          ( DownstreamStackBusLane[6][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane15_strm1_data_valid    ( DownstreamStackBusLane[6][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane16_strm0_ready         ( DownstreamStackBusLane[6][16].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane16_strm0_cntl          ( DownstreamStackBusLane[6][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane16_strm0_data          ( DownstreamStackBusLane[6][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane16_strm0_data_valid    ( DownstreamStackBusLane[6][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane16_strm1_ready         ( DownstreamStackBusLane[6][16].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane16_strm1_cntl          ( DownstreamStackBusLane[6][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane16_strm1_data          ( DownstreamStackBusLane[6][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane16_strm1_data_valid    ( DownstreamStackBusLane[6][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane17_strm0_ready         ( DownstreamStackBusLane[6][17].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane17_strm0_cntl          ( DownstreamStackBusLane[6][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane17_strm0_data          ( DownstreamStackBusLane[6][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane17_strm0_data_valid    ( DownstreamStackBusLane[6][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane17_strm1_ready         ( DownstreamStackBusLane[6][17].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane17_strm1_cntl          ( DownstreamStackBusLane[6][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane17_strm1_data          ( DownstreamStackBusLane[6][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane17_strm1_data_valid    ( DownstreamStackBusLane[6][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane18_strm0_ready         ( DownstreamStackBusLane[6][18].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane18_strm0_cntl          ( DownstreamStackBusLane[6][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane18_strm0_data          ( DownstreamStackBusLane[6][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane18_strm0_data_valid    ( DownstreamStackBusLane[6][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane18_strm1_ready         ( DownstreamStackBusLane[6][18].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane18_strm1_cntl          ( DownstreamStackBusLane[6][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane18_strm1_data          ( DownstreamStackBusLane[6][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane18_strm1_data_valid    ( DownstreamStackBusLane[6][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane19_strm0_ready         ( DownstreamStackBusLane[6][19].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane19_strm0_cntl          ( DownstreamStackBusLane[6][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane19_strm0_data          ( DownstreamStackBusLane[6][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane19_strm0_data_valid    ( DownstreamStackBusLane[6][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane19_strm1_ready         ( DownstreamStackBusLane[6][19].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane19_strm1_cntl          ( DownstreamStackBusLane[6][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane19_strm1_data          ( DownstreamStackBusLane[6][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane19_strm1_data_valid    ( DownstreamStackBusLane[6][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane20_strm0_ready         ( DownstreamStackBusLane[6][20].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane20_strm0_cntl          ( DownstreamStackBusLane[6][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane20_strm0_data          ( DownstreamStackBusLane[6][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane20_strm0_data_valid    ( DownstreamStackBusLane[6][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane20_strm1_ready         ( DownstreamStackBusLane[6][20].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane20_strm1_cntl          ( DownstreamStackBusLane[6][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane20_strm1_data          ( DownstreamStackBusLane[6][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane20_strm1_data_valid    ( DownstreamStackBusLane[6][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane21_strm0_ready         ( DownstreamStackBusLane[6][21].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane21_strm0_cntl          ( DownstreamStackBusLane[6][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane21_strm0_data          ( DownstreamStackBusLane[6][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane21_strm0_data_valid    ( DownstreamStackBusLane[6][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane21_strm1_ready         ( DownstreamStackBusLane[6][21].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane21_strm1_cntl          ( DownstreamStackBusLane[6][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane21_strm1_data          ( DownstreamStackBusLane[6][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane21_strm1_data_valid    ( DownstreamStackBusLane[6][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane22_strm0_ready         ( DownstreamStackBusLane[6][22].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane22_strm0_cntl          ( DownstreamStackBusLane[6][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane22_strm0_data          ( DownstreamStackBusLane[6][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane22_strm0_data_valid    ( DownstreamStackBusLane[6][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane22_strm1_ready         ( DownstreamStackBusLane[6][22].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane22_strm1_cntl          ( DownstreamStackBusLane[6][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane22_strm1_data          ( DownstreamStackBusLane[6][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane22_strm1_data_valid    ( DownstreamStackBusLane[6][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane23_strm0_ready         ( DownstreamStackBusLane[6][23].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane23_strm0_cntl          ( DownstreamStackBusLane[6][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane23_strm0_data          ( DownstreamStackBusLane[6][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane23_strm0_data_valid    ( DownstreamStackBusLane[6][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane23_strm1_ready         ( DownstreamStackBusLane[6][23].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane23_strm1_cntl          ( DownstreamStackBusLane[6][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane23_strm1_data          ( DownstreamStackBusLane[6][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane23_strm1_data_valid    ( DownstreamStackBusLane[6][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane24_strm0_ready         ( DownstreamStackBusLane[6][24].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane24_strm0_cntl          ( DownstreamStackBusLane[6][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane24_strm0_data          ( DownstreamStackBusLane[6][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane24_strm0_data_valid    ( DownstreamStackBusLane[6][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane24_strm1_ready         ( DownstreamStackBusLane[6][24].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane24_strm1_cntl          ( DownstreamStackBusLane[6][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane24_strm1_data          ( DownstreamStackBusLane[6][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane24_strm1_data_valid    ( DownstreamStackBusLane[6][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane25_strm0_ready         ( DownstreamStackBusLane[6][25].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane25_strm0_cntl          ( DownstreamStackBusLane[6][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane25_strm0_data          ( DownstreamStackBusLane[6][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane25_strm0_data_valid    ( DownstreamStackBusLane[6][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane25_strm1_ready         ( DownstreamStackBusLane[6][25].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane25_strm1_cntl          ( DownstreamStackBusLane[6][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane25_strm1_data          ( DownstreamStackBusLane[6][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane25_strm1_data_valid    ( DownstreamStackBusLane[6][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane26_strm0_ready         ( DownstreamStackBusLane[6][26].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane26_strm0_cntl          ( DownstreamStackBusLane[6][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane26_strm0_data          ( DownstreamStackBusLane[6][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane26_strm0_data_valid    ( DownstreamStackBusLane[6][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane26_strm1_ready         ( DownstreamStackBusLane[6][26].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane26_strm1_cntl          ( DownstreamStackBusLane[6][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane26_strm1_data          ( DownstreamStackBusLane[6][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane26_strm1_data_valid    ( DownstreamStackBusLane[6][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane27_strm0_ready         ( DownstreamStackBusLane[6][27].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane27_strm0_cntl          ( DownstreamStackBusLane[6][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane27_strm0_data          ( DownstreamStackBusLane[6][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane27_strm0_data_valid    ( DownstreamStackBusLane[6][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane27_strm1_ready         ( DownstreamStackBusLane[6][27].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane27_strm1_cntl          ( DownstreamStackBusLane[6][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane27_strm1_data          ( DownstreamStackBusLane[6][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane27_strm1_data_valid    ( DownstreamStackBusLane[6][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane28_strm0_ready         ( DownstreamStackBusLane[6][28].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane28_strm0_cntl          ( DownstreamStackBusLane[6][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane28_strm0_data          ( DownstreamStackBusLane[6][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane28_strm0_data_valid    ( DownstreamStackBusLane[6][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane28_strm1_ready         ( DownstreamStackBusLane[6][28].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane28_strm1_cntl          ( DownstreamStackBusLane[6][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane28_strm1_data          ( DownstreamStackBusLane[6][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane28_strm1_data_valid    ( DownstreamStackBusLane[6][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane29_strm0_ready         ( DownstreamStackBusLane[6][29].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane29_strm0_cntl          ( DownstreamStackBusLane[6][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane29_strm0_data          ( DownstreamStackBusLane[6][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane29_strm0_data_valid    ( DownstreamStackBusLane[6][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane29_strm1_ready         ( DownstreamStackBusLane[6][29].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane29_strm1_cntl          ( DownstreamStackBusLane[6][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane29_strm1_data          ( DownstreamStackBusLane[6][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane29_strm1_data_valid    ( DownstreamStackBusLane[6][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane30_strm0_ready         ( DownstreamStackBusLane[6][30].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane30_strm0_cntl          ( DownstreamStackBusLane[6][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane30_strm0_data          ( DownstreamStackBusLane[6][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane30_strm0_data_valid    ( DownstreamStackBusLane[6][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane30_strm1_ready         ( DownstreamStackBusLane[6][30].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane30_strm1_cntl          ( DownstreamStackBusLane[6][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane30_strm1_data          ( DownstreamStackBusLane[6][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane30_strm1_data_valid    ( DownstreamStackBusLane[6][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 6, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane31_strm0_ready         ( DownstreamStackBusLane[6][31].pe__std__lane_strm0_ready              ),      
        .std__pe6__lane31_strm0_cntl          ( DownstreamStackBusLane[6][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe6__lane31_strm0_data          ( DownstreamStackBusLane[6][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe6__lane31_strm0_data_valid    ( DownstreamStackBusLane[6][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__std__lane31_strm1_ready         ( DownstreamStackBusLane[6][31].pe__std__lane_strm1_ready              ),      
        .std__pe6__lane31_strm1_cntl          ( DownstreamStackBusLane[6][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe6__lane31_strm1_data          ( DownstreamStackBusLane[6][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe6__lane31_strm1_data_valid    ( DownstreamStackBusLane[6][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane0_strm0_ready         ( DownstreamStackBusLane[7][0].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane0_strm0_cntl          ( DownstreamStackBusLane[7][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane0_strm0_data          ( DownstreamStackBusLane[7][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane0_strm0_data_valid    ( DownstreamStackBusLane[7][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane0_strm1_ready         ( DownstreamStackBusLane[7][0].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane0_strm1_cntl          ( DownstreamStackBusLane[7][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane0_strm1_data          ( DownstreamStackBusLane[7][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane0_strm1_data_valid    ( DownstreamStackBusLane[7][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane1_strm0_ready         ( DownstreamStackBusLane[7][1].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane1_strm0_cntl          ( DownstreamStackBusLane[7][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane1_strm0_data          ( DownstreamStackBusLane[7][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane1_strm0_data_valid    ( DownstreamStackBusLane[7][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane1_strm1_ready         ( DownstreamStackBusLane[7][1].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane1_strm1_cntl          ( DownstreamStackBusLane[7][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane1_strm1_data          ( DownstreamStackBusLane[7][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane1_strm1_data_valid    ( DownstreamStackBusLane[7][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane2_strm0_ready         ( DownstreamStackBusLane[7][2].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane2_strm0_cntl          ( DownstreamStackBusLane[7][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane2_strm0_data          ( DownstreamStackBusLane[7][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane2_strm0_data_valid    ( DownstreamStackBusLane[7][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane2_strm1_ready         ( DownstreamStackBusLane[7][2].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane2_strm1_cntl          ( DownstreamStackBusLane[7][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane2_strm1_data          ( DownstreamStackBusLane[7][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane2_strm1_data_valid    ( DownstreamStackBusLane[7][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane3_strm0_ready         ( DownstreamStackBusLane[7][3].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane3_strm0_cntl          ( DownstreamStackBusLane[7][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane3_strm0_data          ( DownstreamStackBusLane[7][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane3_strm0_data_valid    ( DownstreamStackBusLane[7][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane3_strm1_ready         ( DownstreamStackBusLane[7][3].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane3_strm1_cntl          ( DownstreamStackBusLane[7][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane3_strm1_data          ( DownstreamStackBusLane[7][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane3_strm1_data_valid    ( DownstreamStackBusLane[7][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane4_strm0_ready         ( DownstreamStackBusLane[7][4].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane4_strm0_cntl          ( DownstreamStackBusLane[7][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane4_strm0_data          ( DownstreamStackBusLane[7][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane4_strm0_data_valid    ( DownstreamStackBusLane[7][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane4_strm1_ready         ( DownstreamStackBusLane[7][4].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane4_strm1_cntl          ( DownstreamStackBusLane[7][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane4_strm1_data          ( DownstreamStackBusLane[7][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane4_strm1_data_valid    ( DownstreamStackBusLane[7][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane5_strm0_ready         ( DownstreamStackBusLane[7][5].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane5_strm0_cntl          ( DownstreamStackBusLane[7][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane5_strm0_data          ( DownstreamStackBusLane[7][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane5_strm0_data_valid    ( DownstreamStackBusLane[7][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane5_strm1_ready         ( DownstreamStackBusLane[7][5].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane5_strm1_cntl          ( DownstreamStackBusLane[7][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane5_strm1_data          ( DownstreamStackBusLane[7][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane5_strm1_data_valid    ( DownstreamStackBusLane[7][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane6_strm0_ready         ( DownstreamStackBusLane[7][6].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane6_strm0_cntl          ( DownstreamStackBusLane[7][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane6_strm0_data          ( DownstreamStackBusLane[7][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane6_strm0_data_valid    ( DownstreamStackBusLane[7][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane6_strm1_ready         ( DownstreamStackBusLane[7][6].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane6_strm1_cntl          ( DownstreamStackBusLane[7][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane6_strm1_data          ( DownstreamStackBusLane[7][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane6_strm1_data_valid    ( DownstreamStackBusLane[7][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane7_strm0_ready         ( DownstreamStackBusLane[7][7].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane7_strm0_cntl          ( DownstreamStackBusLane[7][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane7_strm0_data          ( DownstreamStackBusLane[7][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane7_strm0_data_valid    ( DownstreamStackBusLane[7][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane7_strm1_ready         ( DownstreamStackBusLane[7][7].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane7_strm1_cntl          ( DownstreamStackBusLane[7][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane7_strm1_data          ( DownstreamStackBusLane[7][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane7_strm1_data_valid    ( DownstreamStackBusLane[7][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane8_strm0_ready         ( DownstreamStackBusLane[7][8].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane8_strm0_cntl          ( DownstreamStackBusLane[7][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane8_strm0_data          ( DownstreamStackBusLane[7][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane8_strm0_data_valid    ( DownstreamStackBusLane[7][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane8_strm1_ready         ( DownstreamStackBusLane[7][8].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane8_strm1_cntl          ( DownstreamStackBusLane[7][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane8_strm1_data          ( DownstreamStackBusLane[7][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane8_strm1_data_valid    ( DownstreamStackBusLane[7][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane9_strm0_ready         ( DownstreamStackBusLane[7][9].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane9_strm0_cntl          ( DownstreamStackBusLane[7][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane9_strm0_data          ( DownstreamStackBusLane[7][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane9_strm0_data_valid    ( DownstreamStackBusLane[7][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane9_strm1_ready         ( DownstreamStackBusLane[7][9].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane9_strm1_cntl          ( DownstreamStackBusLane[7][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane9_strm1_data          ( DownstreamStackBusLane[7][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane9_strm1_data_valid    ( DownstreamStackBusLane[7][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane10_strm0_ready         ( DownstreamStackBusLane[7][10].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane10_strm0_cntl          ( DownstreamStackBusLane[7][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane10_strm0_data          ( DownstreamStackBusLane[7][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane10_strm0_data_valid    ( DownstreamStackBusLane[7][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane10_strm1_ready         ( DownstreamStackBusLane[7][10].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane10_strm1_cntl          ( DownstreamStackBusLane[7][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane10_strm1_data          ( DownstreamStackBusLane[7][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane10_strm1_data_valid    ( DownstreamStackBusLane[7][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane11_strm0_ready         ( DownstreamStackBusLane[7][11].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane11_strm0_cntl          ( DownstreamStackBusLane[7][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane11_strm0_data          ( DownstreamStackBusLane[7][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane11_strm0_data_valid    ( DownstreamStackBusLane[7][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane11_strm1_ready         ( DownstreamStackBusLane[7][11].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane11_strm1_cntl          ( DownstreamStackBusLane[7][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane11_strm1_data          ( DownstreamStackBusLane[7][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane11_strm1_data_valid    ( DownstreamStackBusLane[7][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane12_strm0_ready         ( DownstreamStackBusLane[7][12].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane12_strm0_cntl          ( DownstreamStackBusLane[7][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane12_strm0_data          ( DownstreamStackBusLane[7][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane12_strm0_data_valid    ( DownstreamStackBusLane[7][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane12_strm1_ready         ( DownstreamStackBusLane[7][12].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane12_strm1_cntl          ( DownstreamStackBusLane[7][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane12_strm1_data          ( DownstreamStackBusLane[7][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane12_strm1_data_valid    ( DownstreamStackBusLane[7][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane13_strm0_ready         ( DownstreamStackBusLane[7][13].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane13_strm0_cntl          ( DownstreamStackBusLane[7][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane13_strm0_data          ( DownstreamStackBusLane[7][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane13_strm0_data_valid    ( DownstreamStackBusLane[7][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane13_strm1_ready         ( DownstreamStackBusLane[7][13].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane13_strm1_cntl          ( DownstreamStackBusLane[7][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane13_strm1_data          ( DownstreamStackBusLane[7][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane13_strm1_data_valid    ( DownstreamStackBusLane[7][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane14_strm0_ready         ( DownstreamStackBusLane[7][14].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane14_strm0_cntl          ( DownstreamStackBusLane[7][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane14_strm0_data          ( DownstreamStackBusLane[7][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane14_strm0_data_valid    ( DownstreamStackBusLane[7][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane14_strm1_ready         ( DownstreamStackBusLane[7][14].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane14_strm1_cntl          ( DownstreamStackBusLane[7][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane14_strm1_data          ( DownstreamStackBusLane[7][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane14_strm1_data_valid    ( DownstreamStackBusLane[7][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane15_strm0_ready         ( DownstreamStackBusLane[7][15].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane15_strm0_cntl          ( DownstreamStackBusLane[7][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane15_strm0_data          ( DownstreamStackBusLane[7][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane15_strm0_data_valid    ( DownstreamStackBusLane[7][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane15_strm1_ready         ( DownstreamStackBusLane[7][15].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane15_strm1_cntl          ( DownstreamStackBusLane[7][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane15_strm1_data          ( DownstreamStackBusLane[7][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane15_strm1_data_valid    ( DownstreamStackBusLane[7][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane16_strm0_ready         ( DownstreamStackBusLane[7][16].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane16_strm0_cntl          ( DownstreamStackBusLane[7][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane16_strm0_data          ( DownstreamStackBusLane[7][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane16_strm0_data_valid    ( DownstreamStackBusLane[7][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane16_strm1_ready         ( DownstreamStackBusLane[7][16].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane16_strm1_cntl          ( DownstreamStackBusLane[7][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane16_strm1_data          ( DownstreamStackBusLane[7][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane16_strm1_data_valid    ( DownstreamStackBusLane[7][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane17_strm0_ready         ( DownstreamStackBusLane[7][17].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane17_strm0_cntl          ( DownstreamStackBusLane[7][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane17_strm0_data          ( DownstreamStackBusLane[7][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane17_strm0_data_valid    ( DownstreamStackBusLane[7][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane17_strm1_ready         ( DownstreamStackBusLane[7][17].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane17_strm1_cntl          ( DownstreamStackBusLane[7][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane17_strm1_data          ( DownstreamStackBusLane[7][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane17_strm1_data_valid    ( DownstreamStackBusLane[7][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane18_strm0_ready         ( DownstreamStackBusLane[7][18].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane18_strm0_cntl          ( DownstreamStackBusLane[7][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane18_strm0_data          ( DownstreamStackBusLane[7][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane18_strm0_data_valid    ( DownstreamStackBusLane[7][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane18_strm1_ready         ( DownstreamStackBusLane[7][18].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane18_strm1_cntl          ( DownstreamStackBusLane[7][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane18_strm1_data          ( DownstreamStackBusLane[7][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane18_strm1_data_valid    ( DownstreamStackBusLane[7][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane19_strm0_ready         ( DownstreamStackBusLane[7][19].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane19_strm0_cntl          ( DownstreamStackBusLane[7][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane19_strm0_data          ( DownstreamStackBusLane[7][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane19_strm0_data_valid    ( DownstreamStackBusLane[7][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane19_strm1_ready         ( DownstreamStackBusLane[7][19].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane19_strm1_cntl          ( DownstreamStackBusLane[7][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane19_strm1_data          ( DownstreamStackBusLane[7][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane19_strm1_data_valid    ( DownstreamStackBusLane[7][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane20_strm0_ready         ( DownstreamStackBusLane[7][20].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane20_strm0_cntl          ( DownstreamStackBusLane[7][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane20_strm0_data          ( DownstreamStackBusLane[7][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane20_strm0_data_valid    ( DownstreamStackBusLane[7][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane20_strm1_ready         ( DownstreamStackBusLane[7][20].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane20_strm1_cntl          ( DownstreamStackBusLane[7][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane20_strm1_data          ( DownstreamStackBusLane[7][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane20_strm1_data_valid    ( DownstreamStackBusLane[7][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane21_strm0_ready         ( DownstreamStackBusLane[7][21].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane21_strm0_cntl          ( DownstreamStackBusLane[7][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane21_strm0_data          ( DownstreamStackBusLane[7][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane21_strm0_data_valid    ( DownstreamStackBusLane[7][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane21_strm1_ready         ( DownstreamStackBusLane[7][21].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane21_strm1_cntl          ( DownstreamStackBusLane[7][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane21_strm1_data          ( DownstreamStackBusLane[7][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane21_strm1_data_valid    ( DownstreamStackBusLane[7][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane22_strm0_ready         ( DownstreamStackBusLane[7][22].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane22_strm0_cntl          ( DownstreamStackBusLane[7][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane22_strm0_data          ( DownstreamStackBusLane[7][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane22_strm0_data_valid    ( DownstreamStackBusLane[7][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane22_strm1_ready         ( DownstreamStackBusLane[7][22].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane22_strm1_cntl          ( DownstreamStackBusLane[7][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane22_strm1_data          ( DownstreamStackBusLane[7][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane22_strm1_data_valid    ( DownstreamStackBusLane[7][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane23_strm0_ready         ( DownstreamStackBusLane[7][23].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane23_strm0_cntl          ( DownstreamStackBusLane[7][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane23_strm0_data          ( DownstreamStackBusLane[7][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane23_strm0_data_valid    ( DownstreamStackBusLane[7][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane23_strm1_ready         ( DownstreamStackBusLane[7][23].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane23_strm1_cntl          ( DownstreamStackBusLane[7][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane23_strm1_data          ( DownstreamStackBusLane[7][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane23_strm1_data_valid    ( DownstreamStackBusLane[7][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane24_strm0_ready         ( DownstreamStackBusLane[7][24].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane24_strm0_cntl          ( DownstreamStackBusLane[7][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane24_strm0_data          ( DownstreamStackBusLane[7][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane24_strm0_data_valid    ( DownstreamStackBusLane[7][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane24_strm1_ready         ( DownstreamStackBusLane[7][24].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane24_strm1_cntl          ( DownstreamStackBusLane[7][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane24_strm1_data          ( DownstreamStackBusLane[7][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane24_strm1_data_valid    ( DownstreamStackBusLane[7][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane25_strm0_ready         ( DownstreamStackBusLane[7][25].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane25_strm0_cntl          ( DownstreamStackBusLane[7][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane25_strm0_data          ( DownstreamStackBusLane[7][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane25_strm0_data_valid    ( DownstreamStackBusLane[7][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane25_strm1_ready         ( DownstreamStackBusLane[7][25].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane25_strm1_cntl          ( DownstreamStackBusLane[7][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane25_strm1_data          ( DownstreamStackBusLane[7][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane25_strm1_data_valid    ( DownstreamStackBusLane[7][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane26_strm0_ready         ( DownstreamStackBusLane[7][26].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane26_strm0_cntl          ( DownstreamStackBusLane[7][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane26_strm0_data          ( DownstreamStackBusLane[7][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane26_strm0_data_valid    ( DownstreamStackBusLane[7][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane26_strm1_ready         ( DownstreamStackBusLane[7][26].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane26_strm1_cntl          ( DownstreamStackBusLane[7][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane26_strm1_data          ( DownstreamStackBusLane[7][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane26_strm1_data_valid    ( DownstreamStackBusLane[7][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane27_strm0_ready         ( DownstreamStackBusLane[7][27].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane27_strm0_cntl          ( DownstreamStackBusLane[7][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane27_strm0_data          ( DownstreamStackBusLane[7][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane27_strm0_data_valid    ( DownstreamStackBusLane[7][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane27_strm1_ready         ( DownstreamStackBusLane[7][27].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane27_strm1_cntl          ( DownstreamStackBusLane[7][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane27_strm1_data          ( DownstreamStackBusLane[7][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane27_strm1_data_valid    ( DownstreamStackBusLane[7][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane28_strm0_ready         ( DownstreamStackBusLane[7][28].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane28_strm0_cntl          ( DownstreamStackBusLane[7][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane28_strm0_data          ( DownstreamStackBusLane[7][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane28_strm0_data_valid    ( DownstreamStackBusLane[7][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane28_strm1_ready         ( DownstreamStackBusLane[7][28].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane28_strm1_cntl          ( DownstreamStackBusLane[7][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane28_strm1_data          ( DownstreamStackBusLane[7][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane28_strm1_data_valid    ( DownstreamStackBusLane[7][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane29_strm0_ready         ( DownstreamStackBusLane[7][29].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane29_strm0_cntl          ( DownstreamStackBusLane[7][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane29_strm0_data          ( DownstreamStackBusLane[7][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane29_strm0_data_valid    ( DownstreamStackBusLane[7][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane29_strm1_ready         ( DownstreamStackBusLane[7][29].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane29_strm1_cntl          ( DownstreamStackBusLane[7][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane29_strm1_data          ( DownstreamStackBusLane[7][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane29_strm1_data_valid    ( DownstreamStackBusLane[7][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane30_strm0_ready         ( DownstreamStackBusLane[7][30].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane30_strm0_cntl          ( DownstreamStackBusLane[7][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane30_strm0_data          ( DownstreamStackBusLane[7][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane30_strm0_data_valid    ( DownstreamStackBusLane[7][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane30_strm1_ready         ( DownstreamStackBusLane[7][30].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane30_strm1_cntl          ( DownstreamStackBusLane[7][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane30_strm1_data          ( DownstreamStackBusLane[7][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane30_strm1_data_valid    ( DownstreamStackBusLane[7][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 7, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane31_strm0_ready         ( DownstreamStackBusLane[7][31].pe__std__lane_strm0_ready              ),      
        .std__pe7__lane31_strm0_cntl          ( DownstreamStackBusLane[7][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe7__lane31_strm0_data          ( DownstreamStackBusLane[7][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe7__lane31_strm0_data_valid    ( DownstreamStackBusLane[7][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__std__lane31_strm1_ready         ( DownstreamStackBusLane[7][31].pe__std__lane_strm1_ready              ),      
        .std__pe7__lane31_strm1_cntl          ( DownstreamStackBusLane[7][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe7__lane31_strm1_data          ( DownstreamStackBusLane[7][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe7__lane31_strm1_data_valid    ( DownstreamStackBusLane[7][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane0_strm0_ready         ( DownstreamStackBusLane[8][0].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane0_strm0_cntl          ( DownstreamStackBusLane[8][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane0_strm0_data          ( DownstreamStackBusLane[8][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane0_strm0_data_valid    ( DownstreamStackBusLane[8][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane0_strm1_ready         ( DownstreamStackBusLane[8][0].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane0_strm1_cntl          ( DownstreamStackBusLane[8][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane0_strm1_data          ( DownstreamStackBusLane[8][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane0_strm1_data_valid    ( DownstreamStackBusLane[8][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane1_strm0_ready         ( DownstreamStackBusLane[8][1].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane1_strm0_cntl          ( DownstreamStackBusLane[8][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane1_strm0_data          ( DownstreamStackBusLane[8][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane1_strm0_data_valid    ( DownstreamStackBusLane[8][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane1_strm1_ready         ( DownstreamStackBusLane[8][1].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane1_strm1_cntl          ( DownstreamStackBusLane[8][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane1_strm1_data          ( DownstreamStackBusLane[8][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane1_strm1_data_valid    ( DownstreamStackBusLane[8][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane2_strm0_ready         ( DownstreamStackBusLane[8][2].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane2_strm0_cntl          ( DownstreamStackBusLane[8][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane2_strm0_data          ( DownstreamStackBusLane[8][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane2_strm0_data_valid    ( DownstreamStackBusLane[8][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane2_strm1_ready         ( DownstreamStackBusLane[8][2].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane2_strm1_cntl          ( DownstreamStackBusLane[8][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane2_strm1_data          ( DownstreamStackBusLane[8][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane2_strm1_data_valid    ( DownstreamStackBusLane[8][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane3_strm0_ready         ( DownstreamStackBusLane[8][3].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane3_strm0_cntl          ( DownstreamStackBusLane[8][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane3_strm0_data          ( DownstreamStackBusLane[8][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane3_strm0_data_valid    ( DownstreamStackBusLane[8][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane3_strm1_ready         ( DownstreamStackBusLane[8][3].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane3_strm1_cntl          ( DownstreamStackBusLane[8][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane3_strm1_data          ( DownstreamStackBusLane[8][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane3_strm1_data_valid    ( DownstreamStackBusLane[8][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane4_strm0_ready         ( DownstreamStackBusLane[8][4].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane4_strm0_cntl          ( DownstreamStackBusLane[8][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane4_strm0_data          ( DownstreamStackBusLane[8][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane4_strm0_data_valid    ( DownstreamStackBusLane[8][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane4_strm1_ready         ( DownstreamStackBusLane[8][4].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane4_strm1_cntl          ( DownstreamStackBusLane[8][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane4_strm1_data          ( DownstreamStackBusLane[8][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane4_strm1_data_valid    ( DownstreamStackBusLane[8][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane5_strm0_ready         ( DownstreamStackBusLane[8][5].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane5_strm0_cntl          ( DownstreamStackBusLane[8][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane5_strm0_data          ( DownstreamStackBusLane[8][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane5_strm0_data_valid    ( DownstreamStackBusLane[8][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane5_strm1_ready         ( DownstreamStackBusLane[8][5].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane5_strm1_cntl          ( DownstreamStackBusLane[8][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane5_strm1_data          ( DownstreamStackBusLane[8][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane5_strm1_data_valid    ( DownstreamStackBusLane[8][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane6_strm0_ready         ( DownstreamStackBusLane[8][6].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane6_strm0_cntl          ( DownstreamStackBusLane[8][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane6_strm0_data          ( DownstreamStackBusLane[8][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane6_strm0_data_valid    ( DownstreamStackBusLane[8][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane6_strm1_ready         ( DownstreamStackBusLane[8][6].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane6_strm1_cntl          ( DownstreamStackBusLane[8][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane6_strm1_data          ( DownstreamStackBusLane[8][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane6_strm1_data_valid    ( DownstreamStackBusLane[8][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane7_strm0_ready         ( DownstreamStackBusLane[8][7].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane7_strm0_cntl          ( DownstreamStackBusLane[8][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane7_strm0_data          ( DownstreamStackBusLane[8][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane7_strm0_data_valid    ( DownstreamStackBusLane[8][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane7_strm1_ready         ( DownstreamStackBusLane[8][7].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane7_strm1_cntl          ( DownstreamStackBusLane[8][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane7_strm1_data          ( DownstreamStackBusLane[8][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane7_strm1_data_valid    ( DownstreamStackBusLane[8][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane8_strm0_ready         ( DownstreamStackBusLane[8][8].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane8_strm0_cntl          ( DownstreamStackBusLane[8][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane8_strm0_data          ( DownstreamStackBusLane[8][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane8_strm0_data_valid    ( DownstreamStackBusLane[8][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane8_strm1_ready         ( DownstreamStackBusLane[8][8].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane8_strm1_cntl          ( DownstreamStackBusLane[8][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane8_strm1_data          ( DownstreamStackBusLane[8][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane8_strm1_data_valid    ( DownstreamStackBusLane[8][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane9_strm0_ready         ( DownstreamStackBusLane[8][9].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane9_strm0_cntl          ( DownstreamStackBusLane[8][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane9_strm0_data          ( DownstreamStackBusLane[8][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane9_strm0_data_valid    ( DownstreamStackBusLane[8][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane9_strm1_ready         ( DownstreamStackBusLane[8][9].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane9_strm1_cntl          ( DownstreamStackBusLane[8][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane9_strm1_data          ( DownstreamStackBusLane[8][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane9_strm1_data_valid    ( DownstreamStackBusLane[8][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane10_strm0_ready         ( DownstreamStackBusLane[8][10].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane10_strm0_cntl          ( DownstreamStackBusLane[8][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane10_strm0_data          ( DownstreamStackBusLane[8][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane10_strm0_data_valid    ( DownstreamStackBusLane[8][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane10_strm1_ready         ( DownstreamStackBusLane[8][10].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane10_strm1_cntl          ( DownstreamStackBusLane[8][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane10_strm1_data          ( DownstreamStackBusLane[8][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane10_strm1_data_valid    ( DownstreamStackBusLane[8][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane11_strm0_ready         ( DownstreamStackBusLane[8][11].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane11_strm0_cntl          ( DownstreamStackBusLane[8][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane11_strm0_data          ( DownstreamStackBusLane[8][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane11_strm0_data_valid    ( DownstreamStackBusLane[8][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane11_strm1_ready         ( DownstreamStackBusLane[8][11].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane11_strm1_cntl          ( DownstreamStackBusLane[8][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane11_strm1_data          ( DownstreamStackBusLane[8][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane11_strm1_data_valid    ( DownstreamStackBusLane[8][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane12_strm0_ready         ( DownstreamStackBusLane[8][12].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane12_strm0_cntl          ( DownstreamStackBusLane[8][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane12_strm0_data          ( DownstreamStackBusLane[8][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane12_strm0_data_valid    ( DownstreamStackBusLane[8][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane12_strm1_ready         ( DownstreamStackBusLane[8][12].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane12_strm1_cntl          ( DownstreamStackBusLane[8][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane12_strm1_data          ( DownstreamStackBusLane[8][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane12_strm1_data_valid    ( DownstreamStackBusLane[8][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane13_strm0_ready         ( DownstreamStackBusLane[8][13].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane13_strm0_cntl          ( DownstreamStackBusLane[8][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane13_strm0_data          ( DownstreamStackBusLane[8][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane13_strm0_data_valid    ( DownstreamStackBusLane[8][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane13_strm1_ready         ( DownstreamStackBusLane[8][13].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane13_strm1_cntl          ( DownstreamStackBusLane[8][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane13_strm1_data          ( DownstreamStackBusLane[8][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane13_strm1_data_valid    ( DownstreamStackBusLane[8][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane14_strm0_ready         ( DownstreamStackBusLane[8][14].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane14_strm0_cntl          ( DownstreamStackBusLane[8][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane14_strm0_data          ( DownstreamStackBusLane[8][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane14_strm0_data_valid    ( DownstreamStackBusLane[8][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane14_strm1_ready         ( DownstreamStackBusLane[8][14].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane14_strm1_cntl          ( DownstreamStackBusLane[8][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane14_strm1_data          ( DownstreamStackBusLane[8][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane14_strm1_data_valid    ( DownstreamStackBusLane[8][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane15_strm0_ready         ( DownstreamStackBusLane[8][15].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane15_strm0_cntl          ( DownstreamStackBusLane[8][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane15_strm0_data          ( DownstreamStackBusLane[8][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane15_strm0_data_valid    ( DownstreamStackBusLane[8][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane15_strm1_ready         ( DownstreamStackBusLane[8][15].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane15_strm1_cntl          ( DownstreamStackBusLane[8][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane15_strm1_data          ( DownstreamStackBusLane[8][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane15_strm1_data_valid    ( DownstreamStackBusLane[8][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane16_strm0_ready         ( DownstreamStackBusLane[8][16].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane16_strm0_cntl          ( DownstreamStackBusLane[8][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane16_strm0_data          ( DownstreamStackBusLane[8][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane16_strm0_data_valid    ( DownstreamStackBusLane[8][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane16_strm1_ready         ( DownstreamStackBusLane[8][16].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane16_strm1_cntl          ( DownstreamStackBusLane[8][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane16_strm1_data          ( DownstreamStackBusLane[8][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane16_strm1_data_valid    ( DownstreamStackBusLane[8][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane17_strm0_ready         ( DownstreamStackBusLane[8][17].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane17_strm0_cntl          ( DownstreamStackBusLane[8][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane17_strm0_data          ( DownstreamStackBusLane[8][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane17_strm0_data_valid    ( DownstreamStackBusLane[8][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane17_strm1_ready         ( DownstreamStackBusLane[8][17].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane17_strm1_cntl          ( DownstreamStackBusLane[8][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane17_strm1_data          ( DownstreamStackBusLane[8][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane17_strm1_data_valid    ( DownstreamStackBusLane[8][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane18_strm0_ready         ( DownstreamStackBusLane[8][18].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane18_strm0_cntl          ( DownstreamStackBusLane[8][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane18_strm0_data          ( DownstreamStackBusLane[8][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane18_strm0_data_valid    ( DownstreamStackBusLane[8][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane18_strm1_ready         ( DownstreamStackBusLane[8][18].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane18_strm1_cntl          ( DownstreamStackBusLane[8][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane18_strm1_data          ( DownstreamStackBusLane[8][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane18_strm1_data_valid    ( DownstreamStackBusLane[8][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane19_strm0_ready         ( DownstreamStackBusLane[8][19].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane19_strm0_cntl          ( DownstreamStackBusLane[8][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane19_strm0_data          ( DownstreamStackBusLane[8][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane19_strm0_data_valid    ( DownstreamStackBusLane[8][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane19_strm1_ready         ( DownstreamStackBusLane[8][19].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane19_strm1_cntl          ( DownstreamStackBusLane[8][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane19_strm1_data          ( DownstreamStackBusLane[8][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane19_strm1_data_valid    ( DownstreamStackBusLane[8][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane20_strm0_ready         ( DownstreamStackBusLane[8][20].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane20_strm0_cntl          ( DownstreamStackBusLane[8][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane20_strm0_data          ( DownstreamStackBusLane[8][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane20_strm0_data_valid    ( DownstreamStackBusLane[8][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane20_strm1_ready         ( DownstreamStackBusLane[8][20].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane20_strm1_cntl          ( DownstreamStackBusLane[8][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane20_strm1_data          ( DownstreamStackBusLane[8][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane20_strm1_data_valid    ( DownstreamStackBusLane[8][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane21_strm0_ready         ( DownstreamStackBusLane[8][21].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane21_strm0_cntl          ( DownstreamStackBusLane[8][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane21_strm0_data          ( DownstreamStackBusLane[8][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane21_strm0_data_valid    ( DownstreamStackBusLane[8][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane21_strm1_ready         ( DownstreamStackBusLane[8][21].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane21_strm1_cntl          ( DownstreamStackBusLane[8][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane21_strm1_data          ( DownstreamStackBusLane[8][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane21_strm1_data_valid    ( DownstreamStackBusLane[8][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane22_strm0_ready         ( DownstreamStackBusLane[8][22].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane22_strm0_cntl          ( DownstreamStackBusLane[8][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane22_strm0_data          ( DownstreamStackBusLane[8][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane22_strm0_data_valid    ( DownstreamStackBusLane[8][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane22_strm1_ready         ( DownstreamStackBusLane[8][22].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane22_strm1_cntl          ( DownstreamStackBusLane[8][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane22_strm1_data          ( DownstreamStackBusLane[8][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane22_strm1_data_valid    ( DownstreamStackBusLane[8][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane23_strm0_ready         ( DownstreamStackBusLane[8][23].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane23_strm0_cntl          ( DownstreamStackBusLane[8][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane23_strm0_data          ( DownstreamStackBusLane[8][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane23_strm0_data_valid    ( DownstreamStackBusLane[8][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane23_strm1_ready         ( DownstreamStackBusLane[8][23].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane23_strm1_cntl          ( DownstreamStackBusLane[8][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane23_strm1_data          ( DownstreamStackBusLane[8][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane23_strm1_data_valid    ( DownstreamStackBusLane[8][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane24_strm0_ready         ( DownstreamStackBusLane[8][24].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane24_strm0_cntl          ( DownstreamStackBusLane[8][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane24_strm0_data          ( DownstreamStackBusLane[8][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane24_strm0_data_valid    ( DownstreamStackBusLane[8][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane24_strm1_ready         ( DownstreamStackBusLane[8][24].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane24_strm1_cntl          ( DownstreamStackBusLane[8][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane24_strm1_data          ( DownstreamStackBusLane[8][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane24_strm1_data_valid    ( DownstreamStackBusLane[8][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane25_strm0_ready         ( DownstreamStackBusLane[8][25].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane25_strm0_cntl          ( DownstreamStackBusLane[8][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane25_strm0_data          ( DownstreamStackBusLane[8][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane25_strm0_data_valid    ( DownstreamStackBusLane[8][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane25_strm1_ready         ( DownstreamStackBusLane[8][25].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane25_strm1_cntl          ( DownstreamStackBusLane[8][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane25_strm1_data          ( DownstreamStackBusLane[8][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane25_strm1_data_valid    ( DownstreamStackBusLane[8][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane26_strm0_ready         ( DownstreamStackBusLane[8][26].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane26_strm0_cntl          ( DownstreamStackBusLane[8][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane26_strm0_data          ( DownstreamStackBusLane[8][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane26_strm0_data_valid    ( DownstreamStackBusLane[8][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane26_strm1_ready         ( DownstreamStackBusLane[8][26].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane26_strm1_cntl          ( DownstreamStackBusLane[8][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane26_strm1_data          ( DownstreamStackBusLane[8][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane26_strm1_data_valid    ( DownstreamStackBusLane[8][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane27_strm0_ready         ( DownstreamStackBusLane[8][27].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane27_strm0_cntl          ( DownstreamStackBusLane[8][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane27_strm0_data          ( DownstreamStackBusLane[8][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane27_strm0_data_valid    ( DownstreamStackBusLane[8][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane27_strm1_ready         ( DownstreamStackBusLane[8][27].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane27_strm1_cntl          ( DownstreamStackBusLane[8][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane27_strm1_data          ( DownstreamStackBusLane[8][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane27_strm1_data_valid    ( DownstreamStackBusLane[8][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane28_strm0_ready         ( DownstreamStackBusLane[8][28].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane28_strm0_cntl          ( DownstreamStackBusLane[8][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane28_strm0_data          ( DownstreamStackBusLane[8][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane28_strm0_data_valid    ( DownstreamStackBusLane[8][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane28_strm1_ready         ( DownstreamStackBusLane[8][28].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane28_strm1_cntl          ( DownstreamStackBusLane[8][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane28_strm1_data          ( DownstreamStackBusLane[8][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane28_strm1_data_valid    ( DownstreamStackBusLane[8][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane29_strm0_ready         ( DownstreamStackBusLane[8][29].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane29_strm0_cntl          ( DownstreamStackBusLane[8][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane29_strm0_data          ( DownstreamStackBusLane[8][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane29_strm0_data_valid    ( DownstreamStackBusLane[8][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane29_strm1_ready         ( DownstreamStackBusLane[8][29].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane29_strm1_cntl          ( DownstreamStackBusLane[8][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane29_strm1_data          ( DownstreamStackBusLane[8][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane29_strm1_data_valid    ( DownstreamStackBusLane[8][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane30_strm0_ready         ( DownstreamStackBusLane[8][30].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane30_strm0_cntl          ( DownstreamStackBusLane[8][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane30_strm0_data          ( DownstreamStackBusLane[8][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane30_strm0_data_valid    ( DownstreamStackBusLane[8][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane30_strm1_ready         ( DownstreamStackBusLane[8][30].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane30_strm1_cntl          ( DownstreamStackBusLane[8][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane30_strm1_data          ( DownstreamStackBusLane[8][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane30_strm1_data_valid    ( DownstreamStackBusLane[8][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 8, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane31_strm0_ready         ( DownstreamStackBusLane[8][31].pe__std__lane_strm0_ready              ),      
        .std__pe8__lane31_strm0_cntl          ( DownstreamStackBusLane[8][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe8__lane31_strm0_data          ( DownstreamStackBusLane[8][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe8__lane31_strm0_data_valid    ( DownstreamStackBusLane[8][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__std__lane31_strm1_ready         ( DownstreamStackBusLane[8][31].pe__std__lane_strm1_ready              ),      
        .std__pe8__lane31_strm1_cntl          ( DownstreamStackBusLane[8][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe8__lane31_strm1_data          ( DownstreamStackBusLane[8][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe8__lane31_strm1_data_valid    ( DownstreamStackBusLane[8][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane0_strm0_ready         ( DownstreamStackBusLane[9][0].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane0_strm0_cntl          ( DownstreamStackBusLane[9][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane0_strm0_data          ( DownstreamStackBusLane[9][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane0_strm0_data_valid    ( DownstreamStackBusLane[9][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane0_strm1_ready         ( DownstreamStackBusLane[9][0].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane0_strm1_cntl          ( DownstreamStackBusLane[9][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane0_strm1_data          ( DownstreamStackBusLane[9][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane0_strm1_data_valid    ( DownstreamStackBusLane[9][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane1_strm0_ready         ( DownstreamStackBusLane[9][1].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane1_strm0_cntl          ( DownstreamStackBusLane[9][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane1_strm0_data          ( DownstreamStackBusLane[9][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane1_strm0_data_valid    ( DownstreamStackBusLane[9][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane1_strm1_ready         ( DownstreamStackBusLane[9][1].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane1_strm1_cntl          ( DownstreamStackBusLane[9][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane1_strm1_data          ( DownstreamStackBusLane[9][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane1_strm1_data_valid    ( DownstreamStackBusLane[9][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane2_strm0_ready         ( DownstreamStackBusLane[9][2].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane2_strm0_cntl          ( DownstreamStackBusLane[9][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane2_strm0_data          ( DownstreamStackBusLane[9][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane2_strm0_data_valid    ( DownstreamStackBusLane[9][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane2_strm1_ready         ( DownstreamStackBusLane[9][2].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane2_strm1_cntl          ( DownstreamStackBusLane[9][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane2_strm1_data          ( DownstreamStackBusLane[9][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane2_strm1_data_valid    ( DownstreamStackBusLane[9][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane3_strm0_ready         ( DownstreamStackBusLane[9][3].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane3_strm0_cntl          ( DownstreamStackBusLane[9][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane3_strm0_data          ( DownstreamStackBusLane[9][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane3_strm0_data_valid    ( DownstreamStackBusLane[9][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane3_strm1_ready         ( DownstreamStackBusLane[9][3].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane3_strm1_cntl          ( DownstreamStackBusLane[9][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane3_strm1_data          ( DownstreamStackBusLane[9][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane3_strm1_data_valid    ( DownstreamStackBusLane[9][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane4_strm0_ready         ( DownstreamStackBusLane[9][4].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane4_strm0_cntl          ( DownstreamStackBusLane[9][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane4_strm0_data          ( DownstreamStackBusLane[9][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane4_strm0_data_valid    ( DownstreamStackBusLane[9][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane4_strm1_ready         ( DownstreamStackBusLane[9][4].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane4_strm1_cntl          ( DownstreamStackBusLane[9][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane4_strm1_data          ( DownstreamStackBusLane[9][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane4_strm1_data_valid    ( DownstreamStackBusLane[9][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane5_strm0_ready         ( DownstreamStackBusLane[9][5].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane5_strm0_cntl          ( DownstreamStackBusLane[9][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane5_strm0_data          ( DownstreamStackBusLane[9][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane5_strm0_data_valid    ( DownstreamStackBusLane[9][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane5_strm1_ready         ( DownstreamStackBusLane[9][5].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane5_strm1_cntl          ( DownstreamStackBusLane[9][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane5_strm1_data          ( DownstreamStackBusLane[9][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane5_strm1_data_valid    ( DownstreamStackBusLane[9][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane6_strm0_ready         ( DownstreamStackBusLane[9][6].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane6_strm0_cntl          ( DownstreamStackBusLane[9][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane6_strm0_data          ( DownstreamStackBusLane[9][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane6_strm0_data_valid    ( DownstreamStackBusLane[9][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane6_strm1_ready         ( DownstreamStackBusLane[9][6].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane6_strm1_cntl          ( DownstreamStackBusLane[9][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane6_strm1_data          ( DownstreamStackBusLane[9][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane6_strm1_data_valid    ( DownstreamStackBusLane[9][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane7_strm0_ready         ( DownstreamStackBusLane[9][7].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane7_strm0_cntl          ( DownstreamStackBusLane[9][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane7_strm0_data          ( DownstreamStackBusLane[9][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane7_strm0_data_valid    ( DownstreamStackBusLane[9][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane7_strm1_ready         ( DownstreamStackBusLane[9][7].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane7_strm1_cntl          ( DownstreamStackBusLane[9][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane7_strm1_data          ( DownstreamStackBusLane[9][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane7_strm1_data_valid    ( DownstreamStackBusLane[9][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane8_strm0_ready         ( DownstreamStackBusLane[9][8].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane8_strm0_cntl          ( DownstreamStackBusLane[9][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane8_strm0_data          ( DownstreamStackBusLane[9][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane8_strm0_data_valid    ( DownstreamStackBusLane[9][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane8_strm1_ready         ( DownstreamStackBusLane[9][8].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane8_strm1_cntl          ( DownstreamStackBusLane[9][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane8_strm1_data          ( DownstreamStackBusLane[9][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane8_strm1_data_valid    ( DownstreamStackBusLane[9][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane9_strm0_ready         ( DownstreamStackBusLane[9][9].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane9_strm0_cntl          ( DownstreamStackBusLane[9][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane9_strm0_data          ( DownstreamStackBusLane[9][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane9_strm0_data_valid    ( DownstreamStackBusLane[9][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane9_strm1_ready         ( DownstreamStackBusLane[9][9].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane9_strm1_cntl          ( DownstreamStackBusLane[9][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane9_strm1_data          ( DownstreamStackBusLane[9][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane9_strm1_data_valid    ( DownstreamStackBusLane[9][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane10_strm0_ready         ( DownstreamStackBusLane[9][10].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane10_strm0_cntl          ( DownstreamStackBusLane[9][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane10_strm0_data          ( DownstreamStackBusLane[9][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane10_strm0_data_valid    ( DownstreamStackBusLane[9][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane10_strm1_ready         ( DownstreamStackBusLane[9][10].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane10_strm1_cntl          ( DownstreamStackBusLane[9][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane10_strm1_data          ( DownstreamStackBusLane[9][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane10_strm1_data_valid    ( DownstreamStackBusLane[9][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane11_strm0_ready         ( DownstreamStackBusLane[9][11].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane11_strm0_cntl          ( DownstreamStackBusLane[9][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane11_strm0_data          ( DownstreamStackBusLane[9][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane11_strm0_data_valid    ( DownstreamStackBusLane[9][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane11_strm1_ready         ( DownstreamStackBusLane[9][11].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane11_strm1_cntl          ( DownstreamStackBusLane[9][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane11_strm1_data          ( DownstreamStackBusLane[9][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane11_strm1_data_valid    ( DownstreamStackBusLane[9][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane12_strm0_ready         ( DownstreamStackBusLane[9][12].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane12_strm0_cntl          ( DownstreamStackBusLane[9][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane12_strm0_data          ( DownstreamStackBusLane[9][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane12_strm0_data_valid    ( DownstreamStackBusLane[9][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane12_strm1_ready         ( DownstreamStackBusLane[9][12].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane12_strm1_cntl          ( DownstreamStackBusLane[9][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane12_strm1_data          ( DownstreamStackBusLane[9][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane12_strm1_data_valid    ( DownstreamStackBusLane[9][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane13_strm0_ready         ( DownstreamStackBusLane[9][13].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane13_strm0_cntl          ( DownstreamStackBusLane[9][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane13_strm0_data          ( DownstreamStackBusLane[9][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane13_strm0_data_valid    ( DownstreamStackBusLane[9][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane13_strm1_ready         ( DownstreamStackBusLane[9][13].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane13_strm1_cntl          ( DownstreamStackBusLane[9][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane13_strm1_data          ( DownstreamStackBusLane[9][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane13_strm1_data_valid    ( DownstreamStackBusLane[9][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane14_strm0_ready         ( DownstreamStackBusLane[9][14].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane14_strm0_cntl          ( DownstreamStackBusLane[9][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane14_strm0_data          ( DownstreamStackBusLane[9][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane14_strm0_data_valid    ( DownstreamStackBusLane[9][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane14_strm1_ready         ( DownstreamStackBusLane[9][14].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane14_strm1_cntl          ( DownstreamStackBusLane[9][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane14_strm1_data          ( DownstreamStackBusLane[9][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane14_strm1_data_valid    ( DownstreamStackBusLane[9][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane15_strm0_ready         ( DownstreamStackBusLane[9][15].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane15_strm0_cntl          ( DownstreamStackBusLane[9][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane15_strm0_data          ( DownstreamStackBusLane[9][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane15_strm0_data_valid    ( DownstreamStackBusLane[9][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane15_strm1_ready         ( DownstreamStackBusLane[9][15].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane15_strm1_cntl          ( DownstreamStackBusLane[9][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane15_strm1_data          ( DownstreamStackBusLane[9][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane15_strm1_data_valid    ( DownstreamStackBusLane[9][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane16_strm0_ready         ( DownstreamStackBusLane[9][16].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane16_strm0_cntl          ( DownstreamStackBusLane[9][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane16_strm0_data          ( DownstreamStackBusLane[9][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane16_strm0_data_valid    ( DownstreamStackBusLane[9][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane16_strm1_ready         ( DownstreamStackBusLane[9][16].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane16_strm1_cntl          ( DownstreamStackBusLane[9][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane16_strm1_data          ( DownstreamStackBusLane[9][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane16_strm1_data_valid    ( DownstreamStackBusLane[9][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane17_strm0_ready         ( DownstreamStackBusLane[9][17].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane17_strm0_cntl          ( DownstreamStackBusLane[9][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane17_strm0_data          ( DownstreamStackBusLane[9][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane17_strm0_data_valid    ( DownstreamStackBusLane[9][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane17_strm1_ready         ( DownstreamStackBusLane[9][17].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane17_strm1_cntl          ( DownstreamStackBusLane[9][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane17_strm1_data          ( DownstreamStackBusLane[9][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane17_strm1_data_valid    ( DownstreamStackBusLane[9][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane18_strm0_ready         ( DownstreamStackBusLane[9][18].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane18_strm0_cntl          ( DownstreamStackBusLane[9][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane18_strm0_data          ( DownstreamStackBusLane[9][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane18_strm0_data_valid    ( DownstreamStackBusLane[9][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane18_strm1_ready         ( DownstreamStackBusLane[9][18].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane18_strm1_cntl          ( DownstreamStackBusLane[9][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane18_strm1_data          ( DownstreamStackBusLane[9][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane18_strm1_data_valid    ( DownstreamStackBusLane[9][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane19_strm0_ready         ( DownstreamStackBusLane[9][19].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane19_strm0_cntl          ( DownstreamStackBusLane[9][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane19_strm0_data          ( DownstreamStackBusLane[9][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane19_strm0_data_valid    ( DownstreamStackBusLane[9][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane19_strm1_ready         ( DownstreamStackBusLane[9][19].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane19_strm1_cntl          ( DownstreamStackBusLane[9][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane19_strm1_data          ( DownstreamStackBusLane[9][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane19_strm1_data_valid    ( DownstreamStackBusLane[9][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane20_strm0_ready         ( DownstreamStackBusLane[9][20].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane20_strm0_cntl          ( DownstreamStackBusLane[9][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane20_strm0_data          ( DownstreamStackBusLane[9][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane20_strm0_data_valid    ( DownstreamStackBusLane[9][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane20_strm1_ready         ( DownstreamStackBusLane[9][20].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane20_strm1_cntl          ( DownstreamStackBusLane[9][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane20_strm1_data          ( DownstreamStackBusLane[9][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane20_strm1_data_valid    ( DownstreamStackBusLane[9][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane21_strm0_ready         ( DownstreamStackBusLane[9][21].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane21_strm0_cntl          ( DownstreamStackBusLane[9][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane21_strm0_data          ( DownstreamStackBusLane[9][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane21_strm0_data_valid    ( DownstreamStackBusLane[9][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane21_strm1_ready         ( DownstreamStackBusLane[9][21].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane21_strm1_cntl          ( DownstreamStackBusLane[9][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane21_strm1_data          ( DownstreamStackBusLane[9][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane21_strm1_data_valid    ( DownstreamStackBusLane[9][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane22_strm0_ready         ( DownstreamStackBusLane[9][22].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane22_strm0_cntl          ( DownstreamStackBusLane[9][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane22_strm0_data          ( DownstreamStackBusLane[9][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane22_strm0_data_valid    ( DownstreamStackBusLane[9][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane22_strm1_ready         ( DownstreamStackBusLane[9][22].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane22_strm1_cntl          ( DownstreamStackBusLane[9][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane22_strm1_data          ( DownstreamStackBusLane[9][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane22_strm1_data_valid    ( DownstreamStackBusLane[9][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane23_strm0_ready         ( DownstreamStackBusLane[9][23].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane23_strm0_cntl          ( DownstreamStackBusLane[9][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane23_strm0_data          ( DownstreamStackBusLane[9][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane23_strm0_data_valid    ( DownstreamStackBusLane[9][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane23_strm1_ready         ( DownstreamStackBusLane[9][23].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane23_strm1_cntl          ( DownstreamStackBusLane[9][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane23_strm1_data          ( DownstreamStackBusLane[9][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane23_strm1_data_valid    ( DownstreamStackBusLane[9][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane24_strm0_ready         ( DownstreamStackBusLane[9][24].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane24_strm0_cntl          ( DownstreamStackBusLane[9][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane24_strm0_data          ( DownstreamStackBusLane[9][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane24_strm0_data_valid    ( DownstreamStackBusLane[9][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane24_strm1_ready         ( DownstreamStackBusLane[9][24].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane24_strm1_cntl          ( DownstreamStackBusLane[9][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane24_strm1_data          ( DownstreamStackBusLane[9][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane24_strm1_data_valid    ( DownstreamStackBusLane[9][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane25_strm0_ready         ( DownstreamStackBusLane[9][25].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane25_strm0_cntl          ( DownstreamStackBusLane[9][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane25_strm0_data          ( DownstreamStackBusLane[9][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane25_strm0_data_valid    ( DownstreamStackBusLane[9][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane25_strm1_ready         ( DownstreamStackBusLane[9][25].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane25_strm1_cntl          ( DownstreamStackBusLane[9][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane25_strm1_data          ( DownstreamStackBusLane[9][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane25_strm1_data_valid    ( DownstreamStackBusLane[9][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane26_strm0_ready         ( DownstreamStackBusLane[9][26].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane26_strm0_cntl          ( DownstreamStackBusLane[9][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane26_strm0_data          ( DownstreamStackBusLane[9][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane26_strm0_data_valid    ( DownstreamStackBusLane[9][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane26_strm1_ready         ( DownstreamStackBusLane[9][26].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane26_strm1_cntl          ( DownstreamStackBusLane[9][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane26_strm1_data          ( DownstreamStackBusLane[9][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane26_strm1_data_valid    ( DownstreamStackBusLane[9][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane27_strm0_ready         ( DownstreamStackBusLane[9][27].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane27_strm0_cntl          ( DownstreamStackBusLane[9][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane27_strm0_data          ( DownstreamStackBusLane[9][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane27_strm0_data_valid    ( DownstreamStackBusLane[9][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane27_strm1_ready         ( DownstreamStackBusLane[9][27].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane27_strm1_cntl          ( DownstreamStackBusLane[9][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane27_strm1_data          ( DownstreamStackBusLane[9][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane27_strm1_data_valid    ( DownstreamStackBusLane[9][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane28_strm0_ready         ( DownstreamStackBusLane[9][28].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane28_strm0_cntl          ( DownstreamStackBusLane[9][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane28_strm0_data          ( DownstreamStackBusLane[9][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane28_strm0_data_valid    ( DownstreamStackBusLane[9][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane28_strm1_ready         ( DownstreamStackBusLane[9][28].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane28_strm1_cntl          ( DownstreamStackBusLane[9][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane28_strm1_data          ( DownstreamStackBusLane[9][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane28_strm1_data_valid    ( DownstreamStackBusLane[9][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane29_strm0_ready         ( DownstreamStackBusLane[9][29].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane29_strm0_cntl          ( DownstreamStackBusLane[9][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane29_strm0_data          ( DownstreamStackBusLane[9][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane29_strm0_data_valid    ( DownstreamStackBusLane[9][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane29_strm1_ready         ( DownstreamStackBusLane[9][29].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane29_strm1_cntl          ( DownstreamStackBusLane[9][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane29_strm1_data          ( DownstreamStackBusLane[9][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane29_strm1_data_valid    ( DownstreamStackBusLane[9][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane30_strm0_ready         ( DownstreamStackBusLane[9][30].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane30_strm0_cntl          ( DownstreamStackBusLane[9][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane30_strm0_data          ( DownstreamStackBusLane[9][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane30_strm0_data_valid    ( DownstreamStackBusLane[9][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane30_strm1_ready         ( DownstreamStackBusLane[9][30].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane30_strm1_cntl          ( DownstreamStackBusLane[9][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane30_strm1_data          ( DownstreamStackBusLane[9][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane30_strm1_data_valid    ( DownstreamStackBusLane[9][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 9, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane31_strm0_ready         ( DownstreamStackBusLane[9][31].pe__std__lane_strm0_ready              ),      
        .std__pe9__lane31_strm0_cntl          ( DownstreamStackBusLane[9][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe9__lane31_strm0_data          ( DownstreamStackBusLane[9][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe9__lane31_strm0_data_valid    ( DownstreamStackBusLane[9][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__std__lane31_strm1_ready         ( DownstreamStackBusLane[9][31].pe__std__lane_strm1_ready              ),      
        .std__pe9__lane31_strm1_cntl          ( DownstreamStackBusLane[9][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe9__lane31_strm1_data          ( DownstreamStackBusLane[9][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe9__lane31_strm1_data_valid    ( DownstreamStackBusLane[9][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane0_strm0_ready         ( DownstreamStackBusLane[10][0].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane0_strm0_cntl          ( DownstreamStackBusLane[10][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane0_strm0_data          ( DownstreamStackBusLane[10][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane0_strm0_data_valid    ( DownstreamStackBusLane[10][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane0_strm1_ready         ( DownstreamStackBusLane[10][0].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane0_strm1_cntl          ( DownstreamStackBusLane[10][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane0_strm1_data          ( DownstreamStackBusLane[10][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane0_strm1_data_valid    ( DownstreamStackBusLane[10][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane1_strm0_ready         ( DownstreamStackBusLane[10][1].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane1_strm0_cntl          ( DownstreamStackBusLane[10][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane1_strm0_data          ( DownstreamStackBusLane[10][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane1_strm0_data_valid    ( DownstreamStackBusLane[10][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane1_strm1_ready         ( DownstreamStackBusLane[10][1].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane1_strm1_cntl          ( DownstreamStackBusLane[10][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane1_strm1_data          ( DownstreamStackBusLane[10][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane1_strm1_data_valid    ( DownstreamStackBusLane[10][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane2_strm0_ready         ( DownstreamStackBusLane[10][2].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane2_strm0_cntl          ( DownstreamStackBusLane[10][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane2_strm0_data          ( DownstreamStackBusLane[10][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane2_strm0_data_valid    ( DownstreamStackBusLane[10][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane2_strm1_ready         ( DownstreamStackBusLane[10][2].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane2_strm1_cntl          ( DownstreamStackBusLane[10][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane2_strm1_data          ( DownstreamStackBusLane[10][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane2_strm1_data_valid    ( DownstreamStackBusLane[10][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane3_strm0_ready         ( DownstreamStackBusLane[10][3].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane3_strm0_cntl          ( DownstreamStackBusLane[10][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane3_strm0_data          ( DownstreamStackBusLane[10][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane3_strm0_data_valid    ( DownstreamStackBusLane[10][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane3_strm1_ready         ( DownstreamStackBusLane[10][3].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane3_strm1_cntl          ( DownstreamStackBusLane[10][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane3_strm1_data          ( DownstreamStackBusLane[10][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane3_strm1_data_valid    ( DownstreamStackBusLane[10][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane4_strm0_ready         ( DownstreamStackBusLane[10][4].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane4_strm0_cntl          ( DownstreamStackBusLane[10][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane4_strm0_data          ( DownstreamStackBusLane[10][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane4_strm0_data_valid    ( DownstreamStackBusLane[10][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane4_strm1_ready         ( DownstreamStackBusLane[10][4].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane4_strm1_cntl          ( DownstreamStackBusLane[10][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane4_strm1_data          ( DownstreamStackBusLane[10][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane4_strm1_data_valid    ( DownstreamStackBusLane[10][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane5_strm0_ready         ( DownstreamStackBusLane[10][5].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane5_strm0_cntl          ( DownstreamStackBusLane[10][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane5_strm0_data          ( DownstreamStackBusLane[10][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane5_strm0_data_valid    ( DownstreamStackBusLane[10][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane5_strm1_ready         ( DownstreamStackBusLane[10][5].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane5_strm1_cntl          ( DownstreamStackBusLane[10][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane5_strm1_data          ( DownstreamStackBusLane[10][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane5_strm1_data_valid    ( DownstreamStackBusLane[10][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane6_strm0_ready         ( DownstreamStackBusLane[10][6].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane6_strm0_cntl          ( DownstreamStackBusLane[10][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane6_strm0_data          ( DownstreamStackBusLane[10][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane6_strm0_data_valid    ( DownstreamStackBusLane[10][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane6_strm1_ready         ( DownstreamStackBusLane[10][6].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane6_strm1_cntl          ( DownstreamStackBusLane[10][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane6_strm1_data          ( DownstreamStackBusLane[10][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane6_strm1_data_valid    ( DownstreamStackBusLane[10][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane7_strm0_ready         ( DownstreamStackBusLane[10][7].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane7_strm0_cntl          ( DownstreamStackBusLane[10][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane7_strm0_data          ( DownstreamStackBusLane[10][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane7_strm0_data_valid    ( DownstreamStackBusLane[10][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane7_strm1_ready         ( DownstreamStackBusLane[10][7].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane7_strm1_cntl          ( DownstreamStackBusLane[10][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane7_strm1_data          ( DownstreamStackBusLane[10][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane7_strm1_data_valid    ( DownstreamStackBusLane[10][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane8_strm0_ready         ( DownstreamStackBusLane[10][8].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane8_strm0_cntl          ( DownstreamStackBusLane[10][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane8_strm0_data          ( DownstreamStackBusLane[10][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane8_strm0_data_valid    ( DownstreamStackBusLane[10][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane8_strm1_ready         ( DownstreamStackBusLane[10][8].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane8_strm1_cntl          ( DownstreamStackBusLane[10][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane8_strm1_data          ( DownstreamStackBusLane[10][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane8_strm1_data_valid    ( DownstreamStackBusLane[10][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane9_strm0_ready         ( DownstreamStackBusLane[10][9].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane9_strm0_cntl          ( DownstreamStackBusLane[10][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane9_strm0_data          ( DownstreamStackBusLane[10][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane9_strm0_data_valid    ( DownstreamStackBusLane[10][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane9_strm1_ready         ( DownstreamStackBusLane[10][9].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane9_strm1_cntl          ( DownstreamStackBusLane[10][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane9_strm1_data          ( DownstreamStackBusLane[10][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane9_strm1_data_valid    ( DownstreamStackBusLane[10][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane10_strm0_ready         ( DownstreamStackBusLane[10][10].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane10_strm0_cntl          ( DownstreamStackBusLane[10][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane10_strm0_data          ( DownstreamStackBusLane[10][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane10_strm0_data_valid    ( DownstreamStackBusLane[10][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane10_strm1_ready         ( DownstreamStackBusLane[10][10].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane10_strm1_cntl          ( DownstreamStackBusLane[10][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane10_strm1_data          ( DownstreamStackBusLane[10][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane10_strm1_data_valid    ( DownstreamStackBusLane[10][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane11_strm0_ready         ( DownstreamStackBusLane[10][11].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane11_strm0_cntl          ( DownstreamStackBusLane[10][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane11_strm0_data          ( DownstreamStackBusLane[10][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane11_strm0_data_valid    ( DownstreamStackBusLane[10][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane11_strm1_ready         ( DownstreamStackBusLane[10][11].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane11_strm1_cntl          ( DownstreamStackBusLane[10][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane11_strm1_data          ( DownstreamStackBusLane[10][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane11_strm1_data_valid    ( DownstreamStackBusLane[10][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane12_strm0_ready         ( DownstreamStackBusLane[10][12].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane12_strm0_cntl          ( DownstreamStackBusLane[10][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane12_strm0_data          ( DownstreamStackBusLane[10][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane12_strm0_data_valid    ( DownstreamStackBusLane[10][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane12_strm1_ready         ( DownstreamStackBusLane[10][12].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane12_strm1_cntl          ( DownstreamStackBusLane[10][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane12_strm1_data          ( DownstreamStackBusLane[10][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane12_strm1_data_valid    ( DownstreamStackBusLane[10][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane13_strm0_ready         ( DownstreamStackBusLane[10][13].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane13_strm0_cntl          ( DownstreamStackBusLane[10][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane13_strm0_data          ( DownstreamStackBusLane[10][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane13_strm0_data_valid    ( DownstreamStackBusLane[10][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane13_strm1_ready         ( DownstreamStackBusLane[10][13].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane13_strm1_cntl          ( DownstreamStackBusLane[10][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane13_strm1_data          ( DownstreamStackBusLane[10][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane13_strm1_data_valid    ( DownstreamStackBusLane[10][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane14_strm0_ready         ( DownstreamStackBusLane[10][14].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane14_strm0_cntl          ( DownstreamStackBusLane[10][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane14_strm0_data          ( DownstreamStackBusLane[10][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane14_strm0_data_valid    ( DownstreamStackBusLane[10][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane14_strm1_ready         ( DownstreamStackBusLane[10][14].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane14_strm1_cntl          ( DownstreamStackBusLane[10][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane14_strm1_data          ( DownstreamStackBusLane[10][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane14_strm1_data_valid    ( DownstreamStackBusLane[10][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane15_strm0_ready         ( DownstreamStackBusLane[10][15].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane15_strm0_cntl          ( DownstreamStackBusLane[10][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane15_strm0_data          ( DownstreamStackBusLane[10][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane15_strm0_data_valid    ( DownstreamStackBusLane[10][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane15_strm1_ready         ( DownstreamStackBusLane[10][15].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane15_strm1_cntl          ( DownstreamStackBusLane[10][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane15_strm1_data          ( DownstreamStackBusLane[10][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane15_strm1_data_valid    ( DownstreamStackBusLane[10][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane16_strm0_ready         ( DownstreamStackBusLane[10][16].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane16_strm0_cntl          ( DownstreamStackBusLane[10][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane16_strm0_data          ( DownstreamStackBusLane[10][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane16_strm0_data_valid    ( DownstreamStackBusLane[10][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane16_strm1_ready         ( DownstreamStackBusLane[10][16].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane16_strm1_cntl          ( DownstreamStackBusLane[10][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane16_strm1_data          ( DownstreamStackBusLane[10][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane16_strm1_data_valid    ( DownstreamStackBusLane[10][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane17_strm0_ready         ( DownstreamStackBusLane[10][17].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane17_strm0_cntl          ( DownstreamStackBusLane[10][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane17_strm0_data          ( DownstreamStackBusLane[10][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane17_strm0_data_valid    ( DownstreamStackBusLane[10][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane17_strm1_ready         ( DownstreamStackBusLane[10][17].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane17_strm1_cntl          ( DownstreamStackBusLane[10][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane17_strm1_data          ( DownstreamStackBusLane[10][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane17_strm1_data_valid    ( DownstreamStackBusLane[10][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane18_strm0_ready         ( DownstreamStackBusLane[10][18].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane18_strm0_cntl          ( DownstreamStackBusLane[10][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane18_strm0_data          ( DownstreamStackBusLane[10][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane18_strm0_data_valid    ( DownstreamStackBusLane[10][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane18_strm1_ready         ( DownstreamStackBusLane[10][18].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane18_strm1_cntl          ( DownstreamStackBusLane[10][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane18_strm1_data          ( DownstreamStackBusLane[10][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane18_strm1_data_valid    ( DownstreamStackBusLane[10][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane19_strm0_ready         ( DownstreamStackBusLane[10][19].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane19_strm0_cntl          ( DownstreamStackBusLane[10][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane19_strm0_data          ( DownstreamStackBusLane[10][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane19_strm0_data_valid    ( DownstreamStackBusLane[10][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane19_strm1_ready         ( DownstreamStackBusLane[10][19].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane19_strm1_cntl          ( DownstreamStackBusLane[10][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane19_strm1_data          ( DownstreamStackBusLane[10][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane19_strm1_data_valid    ( DownstreamStackBusLane[10][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane20_strm0_ready         ( DownstreamStackBusLane[10][20].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane20_strm0_cntl          ( DownstreamStackBusLane[10][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane20_strm0_data          ( DownstreamStackBusLane[10][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane20_strm0_data_valid    ( DownstreamStackBusLane[10][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane20_strm1_ready         ( DownstreamStackBusLane[10][20].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane20_strm1_cntl          ( DownstreamStackBusLane[10][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane20_strm1_data          ( DownstreamStackBusLane[10][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane20_strm1_data_valid    ( DownstreamStackBusLane[10][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane21_strm0_ready         ( DownstreamStackBusLane[10][21].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane21_strm0_cntl          ( DownstreamStackBusLane[10][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane21_strm0_data          ( DownstreamStackBusLane[10][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane21_strm0_data_valid    ( DownstreamStackBusLane[10][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane21_strm1_ready         ( DownstreamStackBusLane[10][21].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane21_strm1_cntl          ( DownstreamStackBusLane[10][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane21_strm1_data          ( DownstreamStackBusLane[10][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane21_strm1_data_valid    ( DownstreamStackBusLane[10][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane22_strm0_ready         ( DownstreamStackBusLane[10][22].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane22_strm0_cntl          ( DownstreamStackBusLane[10][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane22_strm0_data          ( DownstreamStackBusLane[10][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane22_strm0_data_valid    ( DownstreamStackBusLane[10][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane22_strm1_ready         ( DownstreamStackBusLane[10][22].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane22_strm1_cntl          ( DownstreamStackBusLane[10][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane22_strm1_data          ( DownstreamStackBusLane[10][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane22_strm1_data_valid    ( DownstreamStackBusLane[10][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane23_strm0_ready         ( DownstreamStackBusLane[10][23].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane23_strm0_cntl          ( DownstreamStackBusLane[10][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane23_strm0_data          ( DownstreamStackBusLane[10][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane23_strm0_data_valid    ( DownstreamStackBusLane[10][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane23_strm1_ready         ( DownstreamStackBusLane[10][23].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane23_strm1_cntl          ( DownstreamStackBusLane[10][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane23_strm1_data          ( DownstreamStackBusLane[10][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane23_strm1_data_valid    ( DownstreamStackBusLane[10][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane24_strm0_ready         ( DownstreamStackBusLane[10][24].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane24_strm0_cntl          ( DownstreamStackBusLane[10][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane24_strm0_data          ( DownstreamStackBusLane[10][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane24_strm0_data_valid    ( DownstreamStackBusLane[10][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane24_strm1_ready         ( DownstreamStackBusLane[10][24].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane24_strm1_cntl          ( DownstreamStackBusLane[10][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane24_strm1_data          ( DownstreamStackBusLane[10][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane24_strm1_data_valid    ( DownstreamStackBusLane[10][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane25_strm0_ready         ( DownstreamStackBusLane[10][25].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane25_strm0_cntl          ( DownstreamStackBusLane[10][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane25_strm0_data          ( DownstreamStackBusLane[10][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane25_strm0_data_valid    ( DownstreamStackBusLane[10][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane25_strm1_ready         ( DownstreamStackBusLane[10][25].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane25_strm1_cntl          ( DownstreamStackBusLane[10][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane25_strm1_data          ( DownstreamStackBusLane[10][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane25_strm1_data_valid    ( DownstreamStackBusLane[10][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane26_strm0_ready         ( DownstreamStackBusLane[10][26].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane26_strm0_cntl          ( DownstreamStackBusLane[10][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane26_strm0_data          ( DownstreamStackBusLane[10][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane26_strm0_data_valid    ( DownstreamStackBusLane[10][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane26_strm1_ready         ( DownstreamStackBusLane[10][26].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane26_strm1_cntl          ( DownstreamStackBusLane[10][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane26_strm1_data          ( DownstreamStackBusLane[10][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane26_strm1_data_valid    ( DownstreamStackBusLane[10][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane27_strm0_ready         ( DownstreamStackBusLane[10][27].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane27_strm0_cntl          ( DownstreamStackBusLane[10][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane27_strm0_data          ( DownstreamStackBusLane[10][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane27_strm0_data_valid    ( DownstreamStackBusLane[10][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane27_strm1_ready         ( DownstreamStackBusLane[10][27].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane27_strm1_cntl          ( DownstreamStackBusLane[10][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane27_strm1_data          ( DownstreamStackBusLane[10][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane27_strm1_data_valid    ( DownstreamStackBusLane[10][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane28_strm0_ready         ( DownstreamStackBusLane[10][28].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane28_strm0_cntl          ( DownstreamStackBusLane[10][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane28_strm0_data          ( DownstreamStackBusLane[10][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane28_strm0_data_valid    ( DownstreamStackBusLane[10][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane28_strm1_ready         ( DownstreamStackBusLane[10][28].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane28_strm1_cntl          ( DownstreamStackBusLane[10][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane28_strm1_data          ( DownstreamStackBusLane[10][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane28_strm1_data_valid    ( DownstreamStackBusLane[10][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane29_strm0_ready         ( DownstreamStackBusLane[10][29].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane29_strm0_cntl          ( DownstreamStackBusLane[10][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane29_strm0_data          ( DownstreamStackBusLane[10][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane29_strm0_data_valid    ( DownstreamStackBusLane[10][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane29_strm1_ready         ( DownstreamStackBusLane[10][29].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane29_strm1_cntl          ( DownstreamStackBusLane[10][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane29_strm1_data          ( DownstreamStackBusLane[10][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane29_strm1_data_valid    ( DownstreamStackBusLane[10][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane30_strm0_ready         ( DownstreamStackBusLane[10][30].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane30_strm0_cntl          ( DownstreamStackBusLane[10][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane30_strm0_data          ( DownstreamStackBusLane[10][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane30_strm0_data_valid    ( DownstreamStackBusLane[10][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane30_strm1_ready         ( DownstreamStackBusLane[10][30].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane30_strm1_cntl          ( DownstreamStackBusLane[10][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane30_strm1_data          ( DownstreamStackBusLane[10][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane30_strm1_data_valid    ( DownstreamStackBusLane[10][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 10, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane31_strm0_ready         ( DownstreamStackBusLane[10][31].pe__std__lane_strm0_ready              ),      
        .std__pe10__lane31_strm0_cntl          ( DownstreamStackBusLane[10][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe10__lane31_strm0_data          ( DownstreamStackBusLane[10][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe10__lane31_strm0_data_valid    ( DownstreamStackBusLane[10][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__std__lane31_strm1_ready         ( DownstreamStackBusLane[10][31].pe__std__lane_strm1_ready              ),      
        .std__pe10__lane31_strm1_cntl          ( DownstreamStackBusLane[10][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe10__lane31_strm1_data          ( DownstreamStackBusLane[10][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe10__lane31_strm1_data_valid    ( DownstreamStackBusLane[10][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane0_strm0_ready         ( DownstreamStackBusLane[11][0].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane0_strm0_cntl          ( DownstreamStackBusLane[11][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane0_strm0_data          ( DownstreamStackBusLane[11][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane0_strm0_data_valid    ( DownstreamStackBusLane[11][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane0_strm1_ready         ( DownstreamStackBusLane[11][0].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane0_strm1_cntl          ( DownstreamStackBusLane[11][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane0_strm1_data          ( DownstreamStackBusLane[11][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane0_strm1_data_valid    ( DownstreamStackBusLane[11][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane1_strm0_ready         ( DownstreamStackBusLane[11][1].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane1_strm0_cntl          ( DownstreamStackBusLane[11][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane1_strm0_data          ( DownstreamStackBusLane[11][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane1_strm0_data_valid    ( DownstreamStackBusLane[11][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane1_strm1_ready         ( DownstreamStackBusLane[11][1].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane1_strm1_cntl          ( DownstreamStackBusLane[11][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane1_strm1_data          ( DownstreamStackBusLane[11][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane1_strm1_data_valid    ( DownstreamStackBusLane[11][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane2_strm0_ready         ( DownstreamStackBusLane[11][2].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane2_strm0_cntl          ( DownstreamStackBusLane[11][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane2_strm0_data          ( DownstreamStackBusLane[11][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane2_strm0_data_valid    ( DownstreamStackBusLane[11][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane2_strm1_ready         ( DownstreamStackBusLane[11][2].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane2_strm1_cntl          ( DownstreamStackBusLane[11][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane2_strm1_data          ( DownstreamStackBusLane[11][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane2_strm1_data_valid    ( DownstreamStackBusLane[11][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane3_strm0_ready         ( DownstreamStackBusLane[11][3].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane3_strm0_cntl          ( DownstreamStackBusLane[11][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane3_strm0_data          ( DownstreamStackBusLane[11][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane3_strm0_data_valid    ( DownstreamStackBusLane[11][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane3_strm1_ready         ( DownstreamStackBusLane[11][3].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane3_strm1_cntl          ( DownstreamStackBusLane[11][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane3_strm1_data          ( DownstreamStackBusLane[11][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane3_strm1_data_valid    ( DownstreamStackBusLane[11][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane4_strm0_ready         ( DownstreamStackBusLane[11][4].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane4_strm0_cntl          ( DownstreamStackBusLane[11][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane4_strm0_data          ( DownstreamStackBusLane[11][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane4_strm0_data_valid    ( DownstreamStackBusLane[11][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane4_strm1_ready         ( DownstreamStackBusLane[11][4].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane4_strm1_cntl          ( DownstreamStackBusLane[11][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane4_strm1_data          ( DownstreamStackBusLane[11][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane4_strm1_data_valid    ( DownstreamStackBusLane[11][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane5_strm0_ready         ( DownstreamStackBusLane[11][5].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane5_strm0_cntl          ( DownstreamStackBusLane[11][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane5_strm0_data          ( DownstreamStackBusLane[11][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane5_strm0_data_valid    ( DownstreamStackBusLane[11][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane5_strm1_ready         ( DownstreamStackBusLane[11][5].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane5_strm1_cntl          ( DownstreamStackBusLane[11][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane5_strm1_data          ( DownstreamStackBusLane[11][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane5_strm1_data_valid    ( DownstreamStackBusLane[11][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane6_strm0_ready         ( DownstreamStackBusLane[11][6].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane6_strm0_cntl          ( DownstreamStackBusLane[11][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane6_strm0_data          ( DownstreamStackBusLane[11][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane6_strm0_data_valid    ( DownstreamStackBusLane[11][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane6_strm1_ready         ( DownstreamStackBusLane[11][6].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane6_strm1_cntl          ( DownstreamStackBusLane[11][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane6_strm1_data          ( DownstreamStackBusLane[11][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane6_strm1_data_valid    ( DownstreamStackBusLane[11][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane7_strm0_ready         ( DownstreamStackBusLane[11][7].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane7_strm0_cntl          ( DownstreamStackBusLane[11][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane7_strm0_data          ( DownstreamStackBusLane[11][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane7_strm0_data_valid    ( DownstreamStackBusLane[11][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane7_strm1_ready         ( DownstreamStackBusLane[11][7].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane7_strm1_cntl          ( DownstreamStackBusLane[11][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane7_strm1_data          ( DownstreamStackBusLane[11][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane7_strm1_data_valid    ( DownstreamStackBusLane[11][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane8_strm0_ready         ( DownstreamStackBusLane[11][8].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane8_strm0_cntl          ( DownstreamStackBusLane[11][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane8_strm0_data          ( DownstreamStackBusLane[11][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane8_strm0_data_valid    ( DownstreamStackBusLane[11][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane8_strm1_ready         ( DownstreamStackBusLane[11][8].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane8_strm1_cntl          ( DownstreamStackBusLane[11][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane8_strm1_data          ( DownstreamStackBusLane[11][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane8_strm1_data_valid    ( DownstreamStackBusLane[11][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane9_strm0_ready         ( DownstreamStackBusLane[11][9].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane9_strm0_cntl          ( DownstreamStackBusLane[11][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane9_strm0_data          ( DownstreamStackBusLane[11][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane9_strm0_data_valid    ( DownstreamStackBusLane[11][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane9_strm1_ready         ( DownstreamStackBusLane[11][9].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane9_strm1_cntl          ( DownstreamStackBusLane[11][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane9_strm1_data          ( DownstreamStackBusLane[11][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane9_strm1_data_valid    ( DownstreamStackBusLane[11][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane10_strm0_ready         ( DownstreamStackBusLane[11][10].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane10_strm0_cntl          ( DownstreamStackBusLane[11][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane10_strm0_data          ( DownstreamStackBusLane[11][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane10_strm0_data_valid    ( DownstreamStackBusLane[11][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane10_strm1_ready         ( DownstreamStackBusLane[11][10].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane10_strm1_cntl          ( DownstreamStackBusLane[11][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane10_strm1_data          ( DownstreamStackBusLane[11][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane10_strm1_data_valid    ( DownstreamStackBusLane[11][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane11_strm0_ready         ( DownstreamStackBusLane[11][11].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane11_strm0_cntl          ( DownstreamStackBusLane[11][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane11_strm0_data          ( DownstreamStackBusLane[11][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane11_strm0_data_valid    ( DownstreamStackBusLane[11][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane11_strm1_ready         ( DownstreamStackBusLane[11][11].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane11_strm1_cntl          ( DownstreamStackBusLane[11][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane11_strm1_data          ( DownstreamStackBusLane[11][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane11_strm1_data_valid    ( DownstreamStackBusLane[11][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane12_strm0_ready         ( DownstreamStackBusLane[11][12].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane12_strm0_cntl          ( DownstreamStackBusLane[11][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane12_strm0_data          ( DownstreamStackBusLane[11][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane12_strm0_data_valid    ( DownstreamStackBusLane[11][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane12_strm1_ready         ( DownstreamStackBusLane[11][12].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane12_strm1_cntl          ( DownstreamStackBusLane[11][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane12_strm1_data          ( DownstreamStackBusLane[11][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane12_strm1_data_valid    ( DownstreamStackBusLane[11][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane13_strm0_ready         ( DownstreamStackBusLane[11][13].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane13_strm0_cntl          ( DownstreamStackBusLane[11][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane13_strm0_data          ( DownstreamStackBusLane[11][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane13_strm0_data_valid    ( DownstreamStackBusLane[11][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane13_strm1_ready         ( DownstreamStackBusLane[11][13].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane13_strm1_cntl          ( DownstreamStackBusLane[11][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane13_strm1_data          ( DownstreamStackBusLane[11][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane13_strm1_data_valid    ( DownstreamStackBusLane[11][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane14_strm0_ready         ( DownstreamStackBusLane[11][14].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane14_strm0_cntl          ( DownstreamStackBusLane[11][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane14_strm0_data          ( DownstreamStackBusLane[11][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane14_strm0_data_valid    ( DownstreamStackBusLane[11][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane14_strm1_ready         ( DownstreamStackBusLane[11][14].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane14_strm1_cntl          ( DownstreamStackBusLane[11][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane14_strm1_data          ( DownstreamStackBusLane[11][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane14_strm1_data_valid    ( DownstreamStackBusLane[11][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane15_strm0_ready         ( DownstreamStackBusLane[11][15].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane15_strm0_cntl          ( DownstreamStackBusLane[11][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane15_strm0_data          ( DownstreamStackBusLane[11][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane15_strm0_data_valid    ( DownstreamStackBusLane[11][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane15_strm1_ready         ( DownstreamStackBusLane[11][15].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane15_strm1_cntl          ( DownstreamStackBusLane[11][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane15_strm1_data          ( DownstreamStackBusLane[11][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane15_strm1_data_valid    ( DownstreamStackBusLane[11][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane16_strm0_ready         ( DownstreamStackBusLane[11][16].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane16_strm0_cntl          ( DownstreamStackBusLane[11][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane16_strm0_data          ( DownstreamStackBusLane[11][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane16_strm0_data_valid    ( DownstreamStackBusLane[11][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane16_strm1_ready         ( DownstreamStackBusLane[11][16].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane16_strm1_cntl          ( DownstreamStackBusLane[11][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane16_strm1_data          ( DownstreamStackBusLane[11][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane16_strm1_data_valid    ( DownstreamStackBusLane[11][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane17_strm0_ready         ( DownstreamStackBusLane[11][17].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane17_strm0_cntl          ( DownstreamStackBusLane[11][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane17_strm0_data          ( DownstreamStackBusLane[11][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane17_strm0_data_valid    ( DownstreamStackBusLane[11][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane17_strm1_ready         ( DownstreamStackBusLane[11][17].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane17_strm1_cntl          ( DownstreamStackBusLane[11][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane17_strm1_data          ( DownstreamStackBusLane[11][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane17_strm1_data_valid    ( DownstreamStackBusLane[11][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane18_strm0_ready         ( DownstreamStackBusLane[11][18].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane18_strm0_cntl          ( DownstreamStackBusLane[11][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane18_strm0_data          ( DownstreamStackBusLane[11][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane18_strm0_data_valid    ( DownstreamStackBusLane[11][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane18_strm1_ready         ( DownstreamStackBusLane[11][18].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane18_strm1_cntl          ( DownstreamStackBusLane[11][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane18_strm1_data          ( DownstreamStackBusLane[11][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane18_strm1_data_valid    ( DownstreamStackBusLane[11][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane19_strm0_ready         ( DownstreamStackBusLane[11][19].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane19_strm0_cntl          ( DownstreamStackBusLane[11][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane19_strm0_data          ( DownstreamStackBusLane[11][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane19_strm0_data_valid    ( DownstreamStackBusLane[11][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane19_strm1_ready         ( DownstreamStackBusLane[11][19].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane19_strm1_cntl          ( DownstreamStackBusLane[11][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane19_strm1_data          ( DownstreamStackBusLane[11][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane19_strm1_data_valid    ( DownstreamStackBusLane[11][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane20_strm0_ready         ( DownstreamStackBusLane[11][20].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane20_strm0_cntl          ( DownstreamStackBusLane[11][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane20_strm0_data          ( DownstreamStackBusLane[11][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane20_strm0_data_valid    ( DownstreamStackBusLane[11][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane20_strm1_ready         ( DownstreamStackBusLane[11][20].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane20_strm1_cntl          ( DownstreamStackBusLane[11][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane20_strm1_data          ( DownstreamStackBusLane[11][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane20_strm1_data_valid    ( DownstreamStackBusLane[11][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane21_strm0_ready         ( DownstreamStackBusLane[11][21].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane21_strm0_cntl          ( DownstreamStackBusLane[11][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane21_strm0_data          ( DownstreamStackBusLane[11][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane21_strm0_data_valid    ( DownstreamStackBusLane[11][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane21_strm1_ready         ( DownstreamStackBusLane[11][21].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane21_strm1_cntl          ( DownstreamStackBusLane[11][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane21_strm1_data          ( DownstreamStackBusLane[11][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane21_strm1_data_valid    ( DownstreamStackBusLane[11][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane22_strm0_ready         ( DownstreamStackBusLane[11][22].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane22_strm0_cntl          ( DownstreamStackBusLane[11][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane22_strm0_data          ( DownstreamStackBusLane[11][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane22_strm0_data_valid    ( DownstreamStackBusLane[11][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane22_strm1_ready         ( DownstreamStackBusLane[11][22].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane22_strm1_cntl          ( DownstreamStackBusLane[11][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane22_strm1_data          ( DownstreamStackBusLane[11][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane22_strm1_data_valid    ( DownstreamStackBusLane[11][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane23_strm0_ready         ( DownstreamStackBusLane[11][23].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane23_strm0_cntl          ( DownstreamStackBusLane[11][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane23_strm0_data          ( DownstreamStackBusLane[11][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane23_strm0_data_valid    ( DownstreamStackBusLane[11][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane23_strm1_ready         ( DownstreamStackBusLane[11][23].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane23_strm1_cntl          ( DownstreamStackBusLane[11][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane23_strm1_data          ( DownstreamStackBusLane[11][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane23_strm1_data_valid    ( DownstreamStackBusLane[11][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane24_strm0_ready         ( DownstreamStackBusLane[11][24].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane24_strm0_cntl          ( DownstreamStackBusLane[11][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane24_strm0_data          ( DownstreamStackBusLane[11][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane24_strm0_data_valid    ( DownstreamStackBusLane[11][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane24_strm1_ready         ( DownstreamStackBusLane[11][24].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane24_strm1_cntl          ( DownstreamStackBusLane[11][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane24_strm1_data          ( DownstreamStackBusLane[11][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane24_strm1_data_valid    ( DownstreamStackBusLane[11][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane25_strm0_ready         ( DownstreamStackBusLane[11][25].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane25_strm0_cntl          ( DownstreamStackBusLane[11][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane25_strm0_data          ( DownstreamStackBusLane[11][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane25_strm0_data_valid    ( DownstreamStackBusLane[11][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane25_strm1_ready         ( DownstreamStackBusLane[11][25].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane25_strm1_cntl          ( DownstreamStackBusLane[11][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane25_strm1_data          ( DownstreamStackBusLane[11][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane25_strm1_data_valid    ( DownstreamStackBusLane[11][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane26_strm0_ready         ( DownstreamStackBusLane[11][26].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane26_strm0_cntl          ( DownstreamStackBusLane[11][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane26_strm0_data          ( DownstreamStackBusLane[11][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane26_strm0_data_valid    ( DownstreamStackBusLane[11][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane26_strm1_ready         ( DownstreamStackBusLane[11][26].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane26_strm1_cntl          ( DownstreamStackBusLane[11][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane26_strm1_data          ( DownstreamStackBusLane[11][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane26_strm1_data_valid    ( DownstreamStackBusLane[11][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane27_strm0_ready         ( DownstreamStackBusLane[11][27].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane27_strm0_cntl          ( DownstreamStackBusLane[11][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane27_strm0_data          ( DownstreamStackBusLane[11][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane27_strm0_data_valid    ( DownstreamStackBusLane[11][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane27_strm1_ready         ( DownstreamStackBusLane[11][27].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane27_strm1_cntl          ( DownstreamStackBusLane[11][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane27_strm1_data          ( DownstreamStackBusLane[11][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane27_strm1_data_valid    ( DownstreamStackBusLane[11][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane28_strm0_ready         ( DownstreamStackBusLane[11][28].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane28_strm0_cntl          ( DownstreamStackBusLane[11][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane28_strm0_data          ( DownstreamStackBusLane[11][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane28_strm0_data_valid    ( DownstreamStackBusLane[11][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane28_strm1_ready         ( DownstreamStackBusLane[11][28].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane28_strm1_cntl          ( DownstreamStackBusLane[11][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane28_strm1_data          ( DownstreamStackBusLane[11][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane28_strm1_data_valid    ( DownstreamStackBusLane[11][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane29_strm0_ready         ( DownstreamStackBusLane[11][29].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane29_strm0_cntl          ( DownstreamStackBusLane[11][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane29_strm0_data          ( DownstreamStackBusLane[11][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane29_strm0_data_valid    ( DownstreamStackBusLane[11][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane29_strm1_ready         ( DownstreamStackBusLane[11][29].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane29_strm1_cntl          ( DownstreamStackBusLane[11][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane29_strm1_data          ( DownstreamStackBusLane[11][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane29_strm1_data_valid    ( DownstreamStackBusLane[11][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane30_strm0_ready         ( DownstreamStackBusLane[11][30].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane30_strm0_cntl          ( DownstreamStackBusLane[11][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane30_strm0_data          ( DownstreamStackBusLane[11][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane30_strm0_data_valid    ( DownstreamStackBusLane[11][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane30_strm1_ready         ( DownstreamStackBusLane[11][30].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane30_strm1_cntl          ( DownstreamStackBusLane[11][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane30_strm1_data          ( DownstreamStackBusLane[11][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane30_strm1_data_valid    ( DownstreamStackBusLane[11][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 11, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane31_strm0_ready         ( DownstreamStackBusLane[11][31].pe__std__lane_strm0_ready              ),      
        .std__pe11__lane31_strm0_cntl          ( DownstreamStackBusLane[11][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe11__lane31_strm0_data          ( DownstreamStackBusLane[11][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe11__lane31_strm0_data_valid    ( DownstreamStackBusLane[11][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__std__lane31_strm1_ready         ( DownstreamStackBusLane[11][31].pe__std__lane_strm1_ready              ),      
        .std__pe11__lane31_strm1_cntl          ( DownstreamStackBusLane[11][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe11__lane31_strm1_data          ( DownstreamStackBusLane[11][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe11__lane31_strm1_data_valid    ( DownstreamStackBusLane[11][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane0_strm0_ready         ( DownstreamStackBusLane[12][0].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane0_strm0_cntl          ( DownstreamStackBusLane[12][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane0_strm0_data          ( DownstreamStackBusLane[12][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane0_strm0_data_valid    ( DownstreamStackBusLane[12][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane0_strm1_ready         ( DownstreamStackBusLane[12][0].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane0_strm1_cntl          ( DownstreamStackBusLane[12][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane0_strm1_data          ( DownstreamStackBusLane[12][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane0_strm1_data_valid    ( DownstreamStackBusLane[12][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane1_strm0_ready         ( DownstreamStackBusLane[12][1].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane1_strm0_cntl          ( DownstreamStackBusLane[12][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane1_strm0_data          ( DownstreamStackBusLane[12][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane1_strm0_data_valid    ( DownstreamStackBusLane[12][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane1_strm1_ready         ( DownstreamStackBusLane[12][1].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane1_strm1_cntl          ( DownstreamStackBusLane[12][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane1_strm1_data          ( DownstreamStackBusLane[12][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane1_strm1_data_valid    ( DownstreamStackBusLane[12][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane2_strm0_ready         ( DownstreamStackBusLane[12][2].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane2_strm0_cntl          ( DownstreamStackBusLane[12][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane2_strm0_data          ( DownstreamStackBusLane[12][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane2_strm0_data_valid    ( DownstreamStackBusLane[12][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane2_strm1_ready         ( DownstreamStackBusLane[12][2].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane2_strm1_cntl          ( DownstreamStackBusLane[12][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane2_strm1_data          ( DownstreamStackBusLane[12][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane2_strm1_data_valid    ( DownstreamStackBusLane[12][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane3_strm0_ready         ( DownstreamStackBusLane[12][3].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane3_strm0_cntl          ( DownstreamStackBusLane[12][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane3_strm0_data          ( DownstreamStackBusLane[12][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane3_strm0_data_valid    ( DownstreamStackBusLane[12][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane3_strm1_ready         ( DownstreamStackBusLane[12][3].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane3_strm1_cntl          ( DownstreamStackBusLane[12][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane3_strm1_data          ( DownstreamStackBusLane[12][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane3_strm1_data_valid    ( DownstreamStackBusLane[12][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane4_strm0_ready         ( DownstreamStackBusLane[12][4].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane4_strm0_cntl          ( DownstreamStackBusLane[12][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane4_strm0_data          ( DownstreamStackBusLane[12][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane4_strm0_data_valid    ( DownstreamStackBusLane[12][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane4_strm1_ready         ( DownstreamStackBusLane[12][4].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane4_strm1_cntl          ( DownstreamStackBusLane[12][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane4_strm1_data          ( DownstreamStackBusLane[12][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane4_strm1_data_valid    ( DownstreamStackBusLane[12][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane5_strm0_ready         ( DownstreamStackBusLane[12][5].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane5_strm0_cntl          ( DownstreamStackBusLane[12][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane5_strm0_data          ( DownstreamStackBusLane[12][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane5_strm0_data_valid    ( DownstreamStackBusLane[12][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane5_strm1_ready         ( DownstreamStackBusLane[12][5].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane5_strm1_cntl          ( DownstreamStackBusLane[12][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane5_strm1_data          ( DownstreamStackBusLane[12][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane5_strm1_data_valid    ( DownstreamStackBusLane[12][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane6_strm0_ready         ( DownstreamStackBusLane[12][6].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane6_strm0_cntl          ( DownstreamStackBusLane[12][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane6_strm0_data          ( DownstreamStackBusLane[12][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane6_strm0_data_valid    ( DownstreamStackBusLane[12][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane6_strm1_ready         ( DownstreamStackBusLane[12][6].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane6_strm1_cntl          ( DownstreamStackBusLane[12][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane6_strm1_data          ( DownstreamStackBusLane[12][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane6_strm1_data_valid    ( DownstreamStackBusLane[12][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane7_strm0_ready         ( DownstreamStackBusLane[12][7].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane7_strm0_cntl          ( DownstreamStackBusLane[12][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane7_strm0_data          ( DownstreamStackBusLane[12][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane7_strm0_data_valid    ( DownstreamStackBusLane[12][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane7_strm1_ready         ( DownstreamStackBusLane[12][7].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane7_strm1_cntl          ( DownstreamStackBusLane[12][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane7_strm1_data          ( DownstreamStackBusLane[12][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane7_strm1_data_valid    ( DownstreamStackBusLane[12][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane8_strm0_ready         ( DownstreamStackBusLane[12][8].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane8_strm0_cntl          ( DownstreamStackBusLane[12][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane8_strm0_data          ( DownstreamStackBusLane[12][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane8_strm0_data_valid    ( DownstreamStackBusLane[12][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane8_strm1_ready         ( DownstreamStackBusLane[12][8].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane8_strm1_cntl          ( DownstreamStackBusLane[12][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane8_strm1_data          ( DownstreamStackBusLane[12][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane8_strm1_data_valid    ( DownstreamStackBusLane[12][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane9_strm0_ready         ( DownstreamStackBusLane[12][9].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane9_strm0_cntl          ( DownstreamStackBusLane[12][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane9_strm0_data          ( DownstreamStackBusLane[12][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane9_strm0_data_valid    ( DownstreamStackBusLane[12][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane9_strm1_ready         ( DownstreamStackBusLane[12][9].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane9_strm1_cntl          ( DownstreamStackBusLane[12][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane9_strm1_data          ( DownstreamStackBusLane[12][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane9_strm1_data_valid    ( DownstreamStackBusLane[12][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane10_strm0_ready         ( DownstreamStackBusLane[12][10].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane10_strm0_cntl          ( DownstreamStackBusLane[12][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane10_strm0_data          ( DownstreamStackBusLane[12][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane10_strm0_data_valid    ( DownstreamStackBusLane[12][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane10_strm1_ready         ( DownstreamStackBusLane[12][10].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane10_strm1_cntl          ( DownstreamStackBusLane[12][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane10_strm1_data          ( DownstreamStackBusLane[12][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane10_strm1_data_valid    ( DownstreamStackBusLane[12][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane11_strm0_ready         ( DownstreamStackBusLane[12][11].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane11_strm0_cntl          ( DownstreamStackBusLane[12][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane11_strm0_data          ( DownstreamStackBusLane[12][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane11_strm0_data_valid    ( DownstreamStackBusLane[12][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane11_strm1_ready         ( DownstreamStackBusLane[12][11].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane11_strm1_cntl          ( DownstreamStackBusLane[12][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane11_strm1_data          ( DownstreamStackBusLane[12][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane11_strm1_data_valid    ( DownstreamStackBusLane[12][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane12_strm0_ready         ( DownstreamStackBusLane[12][12].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane12_strm0_cntl          ( DownstreamStackBusLane[12][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane12_strm0_data          ( DownstreamStackBusLane[12][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane12_strm0_data_valid    ( DownstreamStackBusLane[12][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane12_strm1_ready         ( DownstreamStackBusLane[12][12].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane12_strm1_cntl          ( DownstreamStackBusLane[12][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane12_strm1_data          ( DownstreamStackBusLane[12][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane12_strm1_data_valid    ( DownstreamStackBusLane[12][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane13_strm0_ready         ( DownstreamStackBusLane[12][13].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane13_strm0_cntl          ( DownstreamStackBusLane[12][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane13_strm0_data          ( DownstreamStackBusLane[12][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane13_strm0_data_valid    ( DownstreamStackBusLane[12][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane13_strm1_ready         ( DownstreamStackBusLane[12][13].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane13_strm1_cntl          ( DownstreamStackBusLane[12][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane13_strm1_data          ( DownstreamStackBusLane[12][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane13_strm1_data_valid    ( DownstreamStackBusLane[12][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane14_strm0_ready         ( DownstreamStackBusLane[12][14].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane14_strm0_cntl          ( DownstreamStackBusLane[12][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane14_strm0_data          ( DownstreamStackBusLane[12][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane14_strm0_data_valid    ( DownstreamStackBusLane[12][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane14_strm1_ready         ( DownstreamStackBusLane[12][14].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane14_strm1_cntl          ( DownstreamStackBusLane[12][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane14_strm1_data          ( DownstreamStackBusLane[12][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane14_strm1_data_valid    ( DownstreamStackBusLane[12][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane15_strm0_ready         ( DownstreamStackBusLane[12][15].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane15_strm0_cntl          ( DownstreamStackBusLane[12][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane15_strm0_data          ( DownstreamStackBusLane[12][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane15_strm0_data_valid    ( DownstreamStackBusLane[12][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane15_strm1_ready         ( DownstreamStackBusLane[12][15].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane15_strm1_cntl          ( DownstreamStackBusLane[12][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane15_strm1_data          ( DownstreamStackBusLane[12][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane15_strm1_data_valid    ( DownstreamStackBusLane[12][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane16_strm0_ready         ( DownstreamStackBusLane[12][16].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane16_strm0_cntl          ( DownstreamStackBusLane[12][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane16_strm0_data          ( DownstreamStackBusLane[12][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane16_strm0_data_valid    ( DownstreamStackBusLane[12][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane16_strm1_ready         ( DownstreamStackBusLane[12][16].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane16_strm1_cntl          ( DownstreamStackBusLane[12][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane16_strm1_data          ( DownstreamStackBusLane[12][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane16_strm1_data_valid    ( DownstreamStackBusLane[12][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane17_strm0_ready         ( DownstreamStackBusLane[12][17].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane17_strm0_cntl          ( DownstreamStackBusLane[12][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane17_strm0_data          ( DownstreamStackBusLane[12][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane17_strm0_data_valid    ( DownstreamStackBusLane[12][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane17_strm1_ready         ( DownstreamStackBusLane[12][17].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane17_strm1_cntl          ( DownstreamStackBusLane[12][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane17_strm1_data          ( DownstreamStackBusLane[12][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane17_strm1_data_valid    ( DownstreamStackBusLane[12][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane18_strm0_ready         ( DownstreamStackBusLane[12][18].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane18_strm0_cntl          ( DownstreamStackBusLane[12][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane18_strm0_data          ( DownstreamStackBusLane[12][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane18_strm0_data_valid    ( DownstreamStackBusLane[12][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane18_strm1_ready         ( DownstreamStackBusLane[12][18].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane18_strm1_cntl          ( DownstreamStackBusLane[12][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane18_strm1_data          ( DownstreamStackBusLane[12][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane18_strm1_data_valid    ( DownstreamStackBusLane[12][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane19_strm0_ready         ( DownstreamStackBusLane[12][19].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane19_strm0_cntl          ( DownstreamStackBusLane[12][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane19_strm0_data          ( DownstreamStackBusLane[12][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane19_strm0_data_valid    ( DownstreamStackBusLane[12][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane19_strm1_ready         ( DownstreamStackBusLane[12][19].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane19_strm1_cntl          ( DownstreamStackBusLane[12][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane19_strm1_data          ( DownstreamStackBusLane[12][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane19_strm1_data_valid    ( DownstreamStackBusLane[12][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane20_strm0_ready         ( DownstreamStackBusLane[12][20].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane20_strm0_cntl          ( DownstreamStackBusLane[12][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane20_strm0_data          ( DownstreamStackBusLane[12][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane20_strm0_data_valid    ( DownstreamStackBusLane[12][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane20_strm1_ready         ( DownstreamStackBusLane[12][20].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane20_strm1_cntl          ( DownstreamStackBusLane[12][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane20_strm1_data          ( DownstreamStackBusLane[12][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane20_strm1_data_valid    ( DownstreamStackBusLane[12][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane21_strm0_ready         ( DownstreamStackBusLane[12][21].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane21_strm0_cntl          ( DownstreamStackBusLane[12][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane21_strm0_data          ( DownstreamStackBusLane[12][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane21_strm0_data_valid    ( DownstreamStackBusLane[12][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane21_strm1_ready         ( DownstreamStackBusLane[12][21].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane21_strm1_cntl          ( DownstreamStackBusLane[12][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane21_strm1_data          ( DownstreamStackBusLane[12][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane21_strm1_data_valid    ( DownstreamStackBusLane[12][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane22_strm0_ready         ( DownstreamStackBusLane[12][22].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane22_strm0_cntl          ( DownstreamStackBusLane[12][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane22_strm0_data          ( DownstreamStackBusLane[12][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane22_strm0_data_valid    ( DownstreamStackBusLane[12][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane22_strm1_ready         ( DownstreamStackBusLane[12][22].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane22_strm1_cntl          ( DownstreamStackBusLane[12][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane22_strm1_data          ( DownstreamStackBusLane[12][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane22_strm1_data_valid    ( DownstreamStackBusLane[12][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane23_strm0_ready         ( DownstreamStackBusLane[12][23].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane23_strm0_cntl          ( DownstreamStackBusLane[12][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane23_strm0_data          ( DownstreamStackBusLane[12][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane23_strm0_data_valid    ( DownstreamStackBusLane[12][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane23_strm1_ready         ( DownstreamStackBusLane[12][23].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane23_strm1_cntl          ( DownstreamStackBusLane[12][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane23_strm1_data          ( DownstreamStackBusLane[12][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane23_strm1_data_valid    ( DownstreamStackBusLane[12][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane24_strm0_ready         ( DownstreamStackBusLane[12][24].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane24_strm0_cntl          ( DownstreamStackBusLane[12][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane24_strm0_data          ( DownstreamStackBusLane[12][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane24_strm0_data_valid    ( DownstreamStackBusLane[12][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane24_strm1_ready         ( DownstreamStackBusLane[12][24].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane24_strm1_cntl          ( DownstreamStackBusLane[12][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane24_strm1_data          ( DownstreamStackBusLane[12][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane24_strm1_data_valid    ( DownstreamStackBusLane[12][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane25_strm0_ready         ( DownstreamStackBusLane[12][25].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane25_strm0_cntl          ( DownstreamStackBusLane[12][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane25_strm0_data          ( DownstreamStackBusLane[12][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane25_strm0_data_valid    ( DownstreamStackBusLane[12][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane25_strm1_ready         ( DownstreamStackBusLane[12][25].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane25_strm1_cntl          ( DownstreamStackBusLane[12][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane25_strm1_data          ( DownstreamStackBusLane[12][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane25_strm1_data_valid    ( DownstreamStackBusLane[12][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane26_strm0_ready         ( DownstreamStackBusLane[12][26].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane26_strm0_cntl          ( DownstreamStackBusLane[12][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane26_strm0_data          ( DownstreamStackBusLane[12][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane26_strm0_data_valid    ( DownstreamStackBusLane[12][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane26_strm1_ready         ( DownstreamStackBusLane[12][26].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane26_strm1_cntl          ( DownstreamStackBusLane[12][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane26_strm1_data          ( DownstreamStackBusLane[12][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane26_strm1_data_valid    ( DownstreamStackBusLane[12][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane27_strm0_ready         ( DownstreamStackBusLane[12][27].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane27_strm0_cntl          ( DownstreamStackBusLane[12][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane27_strm0_data          ( DownstreamStackBusLane[12][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane27_strm0_data_valid    ( DownstreamStackBusLane[12][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane27_strm1_ready         ( DownstreamStackBusLane[12][27].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane27_strm1_cntl          ( DownstreamStackBusLane[12][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane27_strm1_data          ( DownstreamStackBusLane[12][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane27_strm1_data_valid    ( DownstreamStackBusLane[12][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane28_strm0_ready         ( DownstreamStackBusLane[12][28].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane28_strm0_cntl          ( DownstreamStackBusLane[12][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane28_strm0_data          ( DownstreamStackBusLane[12][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane28_strm0_data_valid    ( DownstreamStackBusLane[12][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane28_strm1_ready         ( DownstreamStackBusLane[12][28].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane28_strm1_cntl          ( DownstreamStackBusLane[12][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane28_strm1_data          ( DownstreamStackBusLane[12][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane28_strm1_data_valid    ( DownstreamStackBusLane[12][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane29_strm0_ready         ( DownstreamStackBusLane[12][29].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane29_strm0_cntl          ( DownstreamStackBusLane[12][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane29_strm0_data          ( DownstreamStackBusLane[12][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane29_strm0_data_valid    ( DownstreamStackBusLane[12][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane29_strm1_ready         ( DownstreamStackBusLane[12][29].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane29_strm1_cntl          ( DownstreamStackBusLane[12][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane29_strm1_data          ( DownstreamStackBusLane[12][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane29_strm1_data_valid    ( DownstreamStackBusLane[12][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane30_strm0_ready         ( DownstreamStackBusLane[12][30].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane30_strm0_cntl          ( DownstreamStackBusLane[12][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane30_strm0_data          ( DownstreamStackBusLane[12][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane30_strm0_data_valid    ( DownstreamStackBusLane[12][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane30_strm1_ready         ( DownstreamStackBusLane[12][30].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane30_strm1_cntl          ( DownstreamStackBusLane[12][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane30_strm1_data          ( DownstreamStackBusLane[12][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane30_strm1_data_valid    ( DownstreamStackBusLane[12][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 12, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane31_strm0_ready         ( DownstreamStackBusLane[12][31].pe__std__lane_strm0_ready              ),      
        .std__pe12__lane31_strm0_cntl          ( DownstreamStackBusLane[12][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe12__lane31_strm0_data          ( DownstreamStackBusLane[12][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe12__lane31_strm0_data_valid    ( DownstreamStackBusLane[12][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__std__lane31_strm1_ready         ( DownstreamStackBusLane[12][31].pe__std__lane_strm1_ready              ),      
        .std__pe12__lane31_strm1_cntl          ( DownstreamStackBusLane[12][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe12__lane31_strm1_data          ( DownstreamStackBusLane[12][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe12__lane31_strm1_data_valid    ( DownstreamStackBusLane[12][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane0_strm0_ready         ( DownstreamStackBusLane[13][0].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane0_strm0_cntl          ( DownstreamStackBusLane[13][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane0_strm0_data          ( DownstreamStackBusLane[13][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane0_strm0_data_valid    ( DownstreamStackBusLane[13][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane0_strm1_ready         ( DownstreamStackBusLane[13][0].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane0_strm1_cntl          ( DownstreamStackBusLane[13][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane0_strm1_data          ( DownstreamStackBusLane[13][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane0_strm1_data_valid    ( DownstreamStackBusLane[13][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane1_strm0_ready         ( DownstreamStackBusLane[13][1].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane1_strm0_cntl          ( DownstreamStackBusLane[13][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane1_strm0_data          ( DownstreamStackBusLane[13][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane1_strm0_data_valid    ( DownstreamStackBusLane[13][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane1_strm1_ready         ( DownstreamStackBusLane[13][1].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane1_strm1_cntl          ( DownstreamStackBusLane[13][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane1_strm1_data          ( DownstreamStackBusLane[13][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane1_strm1_data_valid    ( DownstreamStackBusLane[13][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane2_strm0_ready         ( DownstreamStackBusLane[13][2].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane2_strm0_cntl          ( DownstreamStackBusLane[13][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane2_strm0_data          ( DownstreamStackBusLane[13][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane2_strm0_data_valid    ( DownstreamStackBusLane[13][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane2_strm1_ready         ( DownstreamStackBusLane[13][2].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane2_strm1_cntl          ( DownstreamStackBusLane[13][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane2_strm1_data          ( DownstreamStackBusLane[13][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane2_strm1_data_valid    ( DownstreamStackBusLane[13][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane3_strm0_ready         ( DownstreamStackBusLane[13][3].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane3_strm0_cntl          ( DownstreamStackBusLane[13][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane3_strm0_data          ( DownstreamStackBusLane[13][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane3_strm0_data_valid    ( DownstreamStackBusLane[13][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane3_strm1_ready         ( DownstreamStackBusLane[13][3].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane3_strm1_cntl          ( DownstreamStackBusLane[13][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane3_strm1_data          ( DownstreamStackBusLane[13][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane3_strm1_data_valid    ( DownstreamStackBusLane[13][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane4_strm0_ready         ( DownstreamStackBusLane[13][4].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane4_strm0_cntl          ( DownstreamStackBusLane[13][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane4_strm0_data          ( DownstreamStackBusLane[13][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane4_strm0_data_valid    ( DownstreamStackBusLane[13][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane4_strm1_ready         ( DownstreamStackBusLane[13][4].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane4_strm1_cntl          ( DownstreamStackBusLane[13][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane4_strm1_data          ( DownstreamStackBusLane[13][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane4_strm1_data_valid    ( DownstreamStackBusLane[13][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane5_strm0_ready         ( DownstreamStackBusLane[13][5].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane5_strm0_cntl          ( DownstreamStackBusLane[13][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane5_strm0_data          ( DownstreamStackBusLane[13][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane5_strm0_data_valid    ( DownstreamStackBusLane[13][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane5_strm1_ready         ( DownstreamStackBusLane[13][5].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane5_strm1_cntl          ( DownstreamStackBusLane[13][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane5_strm1_data          ( DownstreamStackBusLane[13][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane5_strm1_data_valid    ( DownstreamStackBusLane[13][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane6_strm0_ready         ( DownstreamStackBusLane[13][6].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane6_strm0_cntl          ( DownstreamStackBusLane[13][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane6_strm0_data          ( DownstreamStackBusLane[13][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane6_strm0_data_valid    ( DownstreamStackBusLane[13][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane6_strm1_ready         ( DownstreamStackBusLane[13][6].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane6_strm1_cntl          ( DownstreamStackBusLane[13][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane6_strm1_data          ( DownstreamStackBusLane[13][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane6_strm1_data_valid    ( DownstreamStackBusLane[13][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane7_strm0_ready         ( DownstreamStackBusLane[13][7].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane7_strm0_cntl          ( DownstreamStackBusLane[13][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane7_strm0_data          ( DownstreamStackBusLane[13][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane7_strm0_data_valid    ( DownstreamStackBusLane[13][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane7_strm1_ready         ( DownstreamStackBusLane[13][7].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane7_strm1_cntl          ( DownstreamStackBusLane[13][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane7_strm1_data          ( DownstreamStackBusLane[13][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane7_strm1_data_valid    ( DownstreamStackBusLane[13][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane8_strm0_ready         ( DownstreamStackBusLane[13][8].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane8_strm0_cntl          ( DownstreamStackBusLane[13][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane8_strm0_data          ( DownstreamStackBusLane[13][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane8_strm0_data_valid    ( DownstreamStackBusLane[13][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane8_strm1_ready         ( DownstreamStackBusLane[13][8].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane8_strm1_cntl          ( DownstreamStackBusLane[13][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane8_strm1_data          ( DownstreamStackBusLane[13][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane8_strm1_data_valid    ( DownstreamStackBusLane[13][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane9_strm0_ready         ( DownstreamStackBusLane[13][9].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane9_strm0_cntl          ( DownstreamStackBusLane[13][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane9_strm0_data          ( DownstreamStackBusLane[13][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane9_strm0_data_valid    ( DownstreamStackBusLane[13][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane9_strm1_ready         ( DownstreamStackBusLane[13][9].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane9_strm1_cntl          ( DownstreamStackBusLane[13][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane9_strm1_data          ( DownstreamStackBusLane[13][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane9_strm1_data_valid    ( DownstreamStackBusLane[13][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane10_strm0_ready         ( DownstreamStackBusLane[13][10].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane10_strm0_cntl          ( DownstreamStackBusLane[13][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane10_strm0_data          ( DownstreamStackBusLane[13][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane10_strm0_data_valid    ( DownstreamStackBusLane[13][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane10_strm1_ready         ( DownstreamStackBusLane[13][10].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane10_strm1_cntl          ( DownstreamStackBusLane[13][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane10_strm1_data          ( DownstreamStackBusLane[13][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane10_strm1_data_valid    ( DownstreamStackBusLane[13][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane11_strm0_ready         ( DownstreamStackBusLane[13][11].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane11_strm0_cntl          ( DownstreamStackBusLane[13][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane11_strm0_data          ( DownstreamStackBusLane[13][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane11_strm0_data_valid    ( DownstreamStackBusLane[13][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane11_strm1_ready         ( DownstreamStackBusLane[13][11].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane11_strm1_cntl          ( DownstreamStackBusLane[13][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane11_strm1_data          ( DownstreamStackBusLane[13][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane11_strm1_data_valid    ( DownstreamStackBusLane[13][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane12_strm0_ready         ( DownstreamStackBusLane[13][12].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane12_strm0_cntl          ( DownstreamStackBusLane[13][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane12_strm0_data          ( DownstreamStackBusLane[13][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane12_strm0_data_valid    ( DownstreamStackBusLane[13][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane12_strm1_ready         ( DownstreamStackBusLane[13][12].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane12_strm1_cntl          ( DownstreamStackBusLane[13][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane12_strm1_data          ( DownstreamStackBusLane[13][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane12_strm1_data_valid    ( DownstreamStackBusLane[13][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane13_strm0_ready         ( DownstreamStackBusLane[13][13].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane13_strm0_cntl          ( DownstreamStackBusLane[13][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane13_strm0_data          ( DownstreamStackBusLane[13][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane13_strm0_data_valid    ( DownstreamStackBusLane[13][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane13_strm1_ready         ( DownstreamStackBusLane[13][13].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane13_strm1_cntl          ( DownstreamStackBusLane[13][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane13_strm1_data          ( DownstreamStackBusLane[13][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane13_strm1_data_valid    ( DownstreamStackBusLane[13][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane14_strm0_ready         ( DownstreamStackBusLane[13][14].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane14_strm0_cntl          ( DownstreamStackBusLane[13][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane14_strm0_data          ( DownstreamStackBusLane[13][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane14_strm0_data_valid    ( DownstreamStackBusLane[13][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane14_strm1_ready         ( DownstreamStackBusLane[13][14].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane14_strm1_cntl          ( DownstreamStackBusLane[13][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane14_strm1_data          ( DownstreamStackBusLane[13][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane14_strm1_data_valid    ( DownstreamStackBusLane[13][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane15_strm0_ready         ( DownstreamStackBusLane[13][15].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane15_strm0_cntl          ( DownstreamStackBusLane[13][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane15_strm0_data          ( DownstreamStackBusLane[13][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane15_strm0_data_valid    ( DownstreamStackBusLane[13][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane15_strm1_ready         ( DownstreamStackBusLane[13][15].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane15_strm1_cntl          ( DownstreamStackBusLane[13][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane15_strm1_data          ( DownstreamStackBusLane[13][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane15_strm1_data_valid    ( DownstreamStackBusLane[13][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane16_strm0_ready         ( DownstreamStackBusLane[13][16].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane16_strm0_cntl          ( DownstreamStackBusLane[13][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane16_strm0_data          ( DownstreamStackBusLane[13][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane16_strm0_data_valid    ( DownstreamStackBusLane[13][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane16_strm1_ready         ( DownstreamStackBusLane[13][16].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane16_strm1_cntl          ( DownstreamStackBusLane[13][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane16_strm1_data          ( DownstreamStackBusLane[13][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane16_strm1_data_valid    ( DownstreamStackBusLane[13][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane17_strm0_ready         ( DownstreamStackBusLane[13][17].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane17_strm0_cntl          ( DownstreamStackBusLane[13][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane17_strm0_data          ( DownstreamStackBusLane[13][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane17_strm0_data_valid    ( DownstreamStackBusLane[13][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane17_strm1_ready         ( DownstreamStackBusLane[13][17].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane17_strm1_cntl          ( DownstreamStackBusLane[13][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane17_strm1_data          ( DownstreamStackBusLane[13][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane17_strm1_data_valid    ( DownstreamStackBusLane[13][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane18_strm0_ready         ( DownstreamStackBusLane[13][18].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane18_strm0_cntl          ( DownstreamStackBusLane[13][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane18_strm0_data          ( DownstreamStackBusLane[13][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane18_strm0_data_valid    ( DownstreamStackBusLane[13][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane18_strm1_ready         ( DownstreamStackBusLane[13][18].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane18_strm1_cntl          ( DownstreamStackBusLane[13][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane18_strm1_data          ( DownstreamStackBusLane[13][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane18_strm1_data_valid    ( DownstreamStackBusLane[13][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane19_strm0_ready         ( DownstreamStackBusLane[13][19].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane19_strm0_cntl          ( DownstreamStackBusLane[13][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane19_strm0_data          ( DownstreamStackBusLane[13][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane19_strm0_data_valid    ( DownstreamStackBusLane[13][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane19_strm1_ready         ( DownstreamStackBusLane[13][19].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane19_strm1_cntl          ( DownstreamStackBusLane[13][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane19_strm1_data          ( DownstreamStackBusLane[13][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane19_strm1_data_valid    ( DownstreamStackBusLane[13][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane20_strm0_ready         ( DownstreamStackBusLane[13][20].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane20_strm0_cntl          ( DownstreamStackBusLane[13][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane20_strm0_data          ( DownstreamStackBusLane[13][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane20_strm0_data_valid    ( DownstreamStackBusLane[13][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane20_strm1_ready         ( DownstreamStackBusLane[13][20].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane20_strm1_cntl          ( DownstreamStackBusLane[13][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane20_strm1_data          ( DownstreamStackBusLane[13][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane20_strm1_data_valid    ( DownstreamStackBusLane[13][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane21_strm0_ready         ( DownstreamStackBusLane[13][21].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane21_strm0_cntl          ( DownstreamStackBusLane[13][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane21_strm0_data          ( DownstreamStackBusLane[13][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane21_strm0_data_valid    ( DownstreamStackBusLane[13][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane21_strm1_ready         ( DownstreamStackBusLane[13][21].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane21_strm1_cntl          ( DownstreamStackBusLane[13][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane21_strm1_data          ( DownstreamStackBusLane[13][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane21_strm1_data_valid    ( DownstreamStackBusLane[13][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane22_strm0_ready         ( DownstreamStackBusLane[13][22].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane22_strm0_cntl          ( DownstreamStackBusLane[13][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane22_strm0_data          ( DownstreamStackBusLane[13][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane22_strm0_data_valid    ( DownstreamStackBusLane[13][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane22_strm1_ready         ( DownstreamStackBusLane[13][22].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane22_strm1_cntl          ( DownstreamStackBusLane[13][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane22_strm1_data          ( DownstreamStackBusLane[13][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane22_strm1_data_valid    ( DownstreamStackBusLane[13][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane23_strm0_ready         ( DownstreamStackBusLane[13][23].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane23_strm0_cntl          ( DownstreamStackBusLane[13][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane23_strm0_data          ( DownstreamStackBusLane[13][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane23_strm0_data_valid    ( DownstreamStackBusLane[13][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane23_strm1_ready         ( DownstreamStackBusLane[13][23].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane23_strm1_cntl          ( DownstreamStackBusLane[13][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane23_strm1_data          ( DownstreamStackBusLane[13][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane23_strm1_data_valid    ( DownstreamStackBusLane[13][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane24_strm0_ready         ( DownstreamStackBusLane[13][24].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane24_strm0_cntl          ( DownstreamStackBusLane[13][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane24_strm0_data          ( DownstreamStackBusLane[13][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane24_strm0_data_valid    ( DownstreamStackBusLane[13][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane24_strm1_ready         ( DownstreamStackBusLane[13][24].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane24_strm1_cntl          ( DownstreamStackBusLane[13][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane24_strm1_data          ( DownstreamStackBusLane[13][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane24_strm1_data_valid    ( DownstreamStackBusLane[13][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane25_strm0_ready         ( DownstreamStackBusLane[13][25].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane25_strm0_cntl          ( DownstreamStackBusLane[13][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane25_strm0_data          ( DownstreamStackBusLane[13][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane25_strm0_data_valid    ( DownstreamStackBusLane[13][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane25_strm1_ready         ( DownstreamStackBusLane[13][25].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane25_strm1_cntl          ( DownstreamStackBusLane[13][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane25_strm1_data          ( DownstreamStackBusLane[13][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane25_strm1_data_valid    ( DownstreamStackBusLane[13][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane26_strm0_ready         ( DownstreamStackBusLane[13][26].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane26_strm0_cntl          ( DownstreamStackBusLane[13][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane26_strm0_data          ( DownstreamStackBusLane[13][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane26_strm0_data_valid    ( DownstreamStackBusLane[13][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane26_strm1_ready         ( DownstreamStackBusLane[13][26].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane26_strm1_cntl          ( DownstreamStackBusLane[13][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane26_strm1_data          ( DownstreamStackBusLane[13][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane26_strm1_data_valid    ( DownstreamStackBusLane[13][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane27_strm0_ready         ( DownstreamStackBusLane[13][27].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane27_strm0_cntl          ( DownstreamStackBusLane[13][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane27_strm0_data          ( DownstreamStackBusLane[13][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane27_strm0_data_valid    ( DownstreamStackBusLane[13][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane27_strm1_ready         ( DownstreamStackBusLane[13][27].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane27_strm1_cntl          ( DownstreamStackBusLane[13][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane27_strm1_data          ( DownstreamStackBusLane[13][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane27_strm1_data_valid    ( DownstreamStackBusLane[13][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane28_strm0_ready         ( DownstreamStackBusLane[13][28].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane28_strm0_cntl          ( DownstreamStackBusLane[13][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane28_strm0_data          ( DownstreamStackBusLane[13][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane28_strm0_data_valid    ( DownstreamStackBusLane[13][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane28_strm1_ready         ( DownstreamStackBusLane[13][28].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane28_strm1_cntl          ( DownstreamStackBusLane[13][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane28_strm1_data          ( DownstreamStackBusLane[13][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane28_strm1_data_valid    ( DownstreamStackBusLane[13][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane29_strm0_ready         ( DownstreamStackBusLane[13][29].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane29_strm0_cntl          ( DownstreamStackBusLane[13][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane29_strm0_data          ( DownstreamStackBusLane[13][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane29_strm0_data_valid    ( DownstreamStackBusLane[13][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane29_strm1_ready         ( DownstreamStackBusLane[13][29].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane29_strm1_cntl          ( DownstreamStackBusLane[13][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane29_strm1_data          ( DownstreamStackBusLane[13][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane29_strm1_data_valid    ( DownstreamStackBusLane[13][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane30_strm0_ready         ( DownstreamStackBusLane[13][30].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane30_strm0_cntl          ( DownstreamStackBusLane[13][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane30_strm0_data          ( DownstreamStackBusLane[13][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane30_strm0_data_valid    ( DownstreamStackBusLane[13][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane30_strm1_ready         ( DownstreamStackBusLane[13][30].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane30_strm1_cntl          ( DownstreamStackBusLane[13][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane30_strm1_data          ( DownstreamStackBusLane[13][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane30_strm1_data_valid    ( DownstreamStackBusLane[13][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 13, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane31_strm0_ready         ( DownstreamStackBusLane[13][31].pe__std__lane_strm0_ready              ),      
        .std__pe13__lane31_strm0_cntl          ( DownstreamStackBusLane[13][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe13__lane31_strm0_data          ( DownstreamStackBusLane[13][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe13__lane31_strm0_data_valid    ( DownstreamStackBusLane[13][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__std__lane31_strm1_ready         ( DownstreamStackBusLane[13][31].pe__std__lane_strm1_ready              ),      
        .std__pe13__lane31_strm1_cntl          ( DownstreamStackBusLane[13][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe13__lane31_strm1_data          ( DownstreamStackBusLane[13][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe13__lane31_strm1_data_valid    ( DownstreamStackBusLane[13][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane0_strm0_ready         ( DownstreamStackBusLane[14][0].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane0_strm0_cntl          ( DownstreamStackBusLane[14][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane0_strm0_data          ( DownstreamStackBusLane[14][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane0_strm0_data_valid    ( DownstreamStackBusLane[14][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane0_strm1_ready         ( DownstreamStackBusLane[14][0].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane0_strm1_cntl          ( DownstreamStackBusLane[14][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane0_strm1_data          ( DownstreamStackBusLane[14][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane0_strm1_data_valid    ( DownstreamStackBusLane[14][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane1_strm0_ready         ( DownstreamStackBusLane[14][1].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane1_strm0_cntl          ( DownstreamStackBusLane[14][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane1_strm0_data          ( DownstreamStackBusLane[14][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane1_strm0_data_valid    ( DownstreamStackBusLane[14][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane1_strm1_ready         ( DownstreamStackBusLane[14][1].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane1_strm1_cntl          ( DownstreamStackBusLane[14][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane1_strm1_data          ( DownstreamStackBusLane[14][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane1_strm1_data_valid    ( DownstreamStackBusLane[14][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane2_strm0_ready         ( DownstreamStackBusLane[14][2].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane2_strm0_cntl          ( DownstreamStackBusLane[14][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane2_strm0_data          ( DownstreamStackBusLane[14][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane2_strm0_data_valid    ( DownstreamStackBusLane[14][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane2_strm1_ready         ( DownstreamStackBusLane[14][2].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane2_strm1_cntl          ( DownstreamStackBusLane[14][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane2_strm1_data          ( DownstreamStackBusLane[14][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane2_strm1_data_valid    ( DownstreamStackBusLane[14][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane3_strm0_ready         ( DownstreamStackBusLane[14][3].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane3_strm0_cntl          ( DownstreamStackBusLane[14][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane3_strm0_data          ( DownstreamStackBusLane[14][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane3_strm0_data_valid    ( DownstreamStackBusLane[14][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane3_strm1_ready         ( DownstreamStackBusLane[14][3].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane3_strm1_cntl          ( DownstreamStackBusLane[14][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane3_strm1_data          ( DownstreamStackBusLane[14][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane3_strm1_data_valid    ( DownstreamStackBusLane[14][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane4_strm0_ready         ( DownstreamStackBusLane[14][4].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane4_strm0_cntl          ( DownstreamStackBusLane[14][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane4_strm0_data          ( DownstreamStackBusLane[14][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane4_strm0_data_valid    ( DownstreamStackBusLane[14][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane4_strm1_ready         ( DownstreamStackBusLane[14][4].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane4_strm1_cntl          ( DownstreamStackBusLane[14][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane4_strm1_data          ( DownstreamStackBusLane[14][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane4_strm1_data_valid    ( DownstreamStackBusLane[14][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane5_strm0_ready         ( DownstreamStackBusLane[14][5].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane5_strm0_cntl          ( DownstreamStackBusLane[14][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane5_strm0_data          ( DownstreamStackBusLane[14][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane5_strm0_data_valid    ( DownstreamStackBusLane[14][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane5_strm1_ready         ( DownstreamStackBusLane[14][5].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane5_strm1_cntl          ( DownstreamStackBusLane[14][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane5_strm1_data          ( DownstreamStackBusLane[14][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane5_strm1_data_valid    ( DownstreamStackBusLane[14][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane6_strm0_ready         ( DownstreamStackBusLane[14][6].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane6_strm0_cntl          ( DownstreamStackBusLane[14][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane6_strm0_data          ( DownstreamStackBusLane[14][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane6_strm0_data_valid    ( DownstreamStackBusLane[14][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane6_strm1_ready         ( DownstreamStackBusLane[14][6].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane6_strm1_cntl          ( DownstreamStackBusLane[14][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane6_strm1_data          ( DownstreamStackBusLane[14][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane6_strm1_data_valid    ( DownstreamStackBusLane[14][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane7_strm0_ready         ( DownstreamStackBusLane[14][7].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane7_strm0_cntl          ( DownstreamStackBusLane[14][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane7_strm0_data          ( DownstreamStackBusLane[14][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane7_strm0_data_valid    ( DownstreamStackBusLane[14][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane7_strm1_ready         ( DownstreamStackBusLane[14][7].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane7_strm1_cntl          ( DownstreamStackBusLane[14][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane7_strm1_data          ( DownstreamStackBusLane[14][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane7_strm1_data_valid    ( DownstreamStackBusLane[14][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane8_strm0_ready         ( DownstreamStackBusLane[14][8].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane8_strm0_cntl          ( DownstreamStackBusLane[14][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane8_strm0_data          ( DownstreamStackBusLane[14][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane8_strm0_data_valid    ( DownstreamStackBusLane[14][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane8_strm1_ready         ( DownstreamStackBusLane[14][8].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane8_strm1_cntl          ( DownstreamStackBusLane[14][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane8_strm1_data          ( DownstreamStackBusLane[14][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane8_strm1_data_valid    ( DownstreamStackBusLane[14][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane9_strm0_ready         ( DownstreamStackBusLane[14][9].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane9_strm0_cntl          ( DownstreamStackBusLane[14][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane9_strm0_data          ( DownstreamStackBusLane[14][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane9_strm0_data_valid    ( DownstreamStackBusLane[14][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane9_strm1_ready         ( DownstreamStackBusLane[14][9].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane9_strm1_cntl          ( DownstreamStackBusLane[14][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane9_strm1_data          ( DownstreamStackBusLane[14][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane9_strm1_data_valid    ( DownstreamStackBusLane[14][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane10_strm0_ready         ( DownstreamStackBusLane[14][10].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane10_strm0_cntl          ( DownstreamStackBusLane[14][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane10_strm0_data          ( DownstreamStackBusLane[14][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane10_strm0_data_valid    ( DownstreamStackBusLane[14][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane10_strm1_ready         ( DownstreamStackBusLane[14][10].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane10_strm1_cntl          ( DownstreamStackBusLane[14][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane10_strm1_data          ( DownstreamStackBusLane[14][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane10_strm1_data_valid    ( DownstreamStackBusLane[14][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane11_strm0_ready         ( DownstreamStackBusLane[14][11].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane11_strm0_cntl          ( DownstreamStackBusLane[14][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane11_strm0_data          ( DownstreamStackBusLane[14][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane11_strm0_data_valid    ( DownstreamStackBusLane[14][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane11_strm1_ready         ( DownstreamStackBusLane[14][11].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane11_strm1_cntl          ( DownstreamStackBusLane[14][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane11_strm1_data          ( DownstreamStackBusLane[14][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane11_strm1_data_valid    ( DownstreamStackBusLane[14][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane12_strm0_ready         ( DownstreamStackBusLane[14][12].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane12_strm0_cntl          ( DownstreamStackBusLane[14][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane12_strm0_data          ( DownstreamStackBusLane[14][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane12_strm0_data_valid    ( DownstreamStackBusLane[14][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane12_strm1_ready         ( DownstreamStackBusLane[14][12].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane12_strm1_cntl          ( DownstreamStackBusLane[14][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane12_strm1_data          ( DownstreamStackBusLane[14][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane12_strm1_data_valid    ( DownstreamStackBusLane[14][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane13_strm0_ready         ( DownstreamStackBusLane[14][13].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane13_strm0_cntl          ( DownstreamStackBusLane[14][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane13_strm0_data          ( DownstreamStackBusLane[14][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane13_strm0_data_valid    ( DownstreamStackBusLane[14][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane13_strm1_ready         ( DownstreamStackBusLane[14][13].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane13_strm1_cntl          ( DownstreamStackBusLane[14][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane13_strm1_data          ( DownstreamStackBusLane[14][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane13_strm1_data_valid    ( DownstreamStackBusLane[14][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane14_strm0_ready         ( DownstreamStackBusLane[14][14].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane14_strm0_cntl          ( DownstreamStackBusLane[14][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane14_strm0_data          ( DownstreamStackBusLane[14][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane14_strm0_data_valid    ( DownstreamStackBusLane[14][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane14_strm1_ready         ( DownstreamStackBusLane[14][14].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane14_strm1_cntl          ( DownstreamStackBusLane[14][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane14_strm1_data          ( DownstreamStackBusLane[14][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane14_strm1_data_valid    ( DownstreamStackBusLane[14][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane15_strm0_ready         ( DownstreamStackBusLane[14][15].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane15_strm0_cntl          ( DownstreamStackBusLane[14][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane15_strm0_data          ( DownstreamStackBusLane[14][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane15_strm0_data_valid    ( DownstreamStackBusLane[14][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane15_strm1_ready         ( DownstreamStackBusLane[14][15].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane15_strm1_cntl          ( DownstreamStackBusLane[14][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane15_strm1_data          ( DownstreamStackBusLane[14][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane15_strm1_data_valid    ( DownstreamStackBusLane[14][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane16_strm0_ready         ( DownstreamStackBusLane[14][16].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane16_strm0_cntl          ( DownstreamStackBusLane[14][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane16_strm0_data          ( DownstreamStackBusLane[14][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane16_strm0_data_valid    ( DownstreamStackBusLane[14][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane16_strm1_ready         ( DownstreamStackBusLane[14][16].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane16_strm1_cntl          ( DownstreamStackBusLane[14][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane16_strm1_data          ( DownstreamStackBusLane[14][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane16_strm1_data_valid    ( DownstreamStackBusLane[14][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane17_strm0_ready         ( DownstreamStackBusLane[14][17].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane17_strm0_cntl          ( DownstreamStackBusLane[14][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane17_strm0_data          ( DownstreamStackBusLane[14][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane17_strm0_data_valid    ( DownstreamStackBusLane[14][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane17_strm1_ready         ( DownstreamStackBusLane[14][17].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane17_strm1_cntl          ( DownstreamStackBusLane[14][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane17_strm1_data          ( DownstreamStackBusLane[14][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane17_strm1_data_valid    ( DownstreamStackBusLane[14][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane18_strm0_ready         ( DownstreamStackBusLane[14][18].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane18_strm0_cntl          ( DownstreamStackBusLane[14][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane18_strm0_data          ( DownstreamStackBusLane[14][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane18_strm0_data_valid    ( DownstreamStackBusLane[14][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane18_strm1_ready         ( DownstreamStackBusLane[14][18].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane18_strm1_cntl          ( DownstreamStackBusLane[14][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane18_strm1_data          ( DownstreamStackBusLane[14][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane18_strm1_data_valid    ( DownstreamStackBusLane[14][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane19_strm0_ready         ( DownstreamStackBusLane[14][19].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane19_strm0_cntl          ( DownstreamStackBusLane[14][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane19_strm0_data          ( DownstreamStackBusLane[14][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane19_strm0_data_valid    ( DownstreamStackBusLane[14][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane19_strm1_ready         ( DownstreamStackBusLane[14][19].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane19_strm1_cntl          ( DownstreamStackBusLane[14][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane19_strm1_data          ( DownstreamStackBusLane[14][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane19_strm1_data_valid    ( DownstreamStackBusLane[14][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane20_strm0_ready         ( DownstreamStackBusLane[14][20].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane20_strm0_cntl          ( DownstreamStackBusLane[14][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane20_strm0_data          ( DownstreamStackBusLane[14][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane20_strm0_data_valid    ( DownstreamStackBusLane[14][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane20_strm1_ready         ( DownstreamStackBusLane[14][20].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane20_strm1_cntl          ( DownstreamStackBusLane[14][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane20_strm1_data          ( DownstreamStackBusLane[14][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane20_strm1_data_valid    ( DownstreamStackBusLane[14][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane21_strm0_ready         ( DownstreamStackBusLane[14][21].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane21_strm0_cntl          ( DownstreamStackBusLane[14][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane21_strm0_data          ( DownstreamStackBusLane[14][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane21_strm0_data_valid    ( DownstreamStackBusLane[14][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane21_strm1_ready         ( DownstreamStackBusLane[14][21].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane21_strm1_cntl          ( DownstreamStackBusLane[14][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane21_strm1_data          ( DownstreamStackBusLane[14][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane21_strm1_data_valid    ( DownstreamStackBusLane[14][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane22_strm0_ready         ( DownstreamStackBusLane[14][22].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane22_strm0_cntl          ( DownstreamStackBusLane[14][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane22_strm0_data          ( DownstreamStackBusLane[14][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane22_strm0_data_valid    ( DownstreamStackBusLane[14][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane22_strm1_ready         ( DownstreamStackBusLane[14][22].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane22_strm1_cntl          ( DownstreamStackBusLane[14][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane22_strm1_data          ( DownstreamStackBusLane[14][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane22_strm1_data_valid    ( DownstreamStackBusLane[14][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane23_strm0_ready         ( DownstreamStackBusLane[14][23].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane23_strm0_cntl          ( DownstreamStackBusLane[14][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane23_strm0_data          ( DownstreamStackBusLane[14][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane23_strm0_data_valid    ( DownstreamStackBusLane[14][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane23_strm1_ready         ( DownstreamStackBusLane[14][23].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane23_strm1_cntl          ( DownstreamStackBusLane[14][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane23_strm1_data          ( DownstreamStackBusLane[14][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane23_strm1_data_valid    ( DownstreamStackBusLane[14][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane24_strm0_ready         ( DownstreamStackBusLane[14][24].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane24_strm0_cntl          ( DownstreamStackBusLane[14][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane24_strm0_data          ( DownstreamStackBusLane[14][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane24_strm0_data_valid    ( DownstreamStackBusLane[14][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane24_strm1_ready         ( DownstreamStackBusLane[14][24].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane24_strm1_cntl          ( DownstreamStackBusLane[14][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane24_strm1_data          ( DownstreamStackBusLane[14][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane24_strm1_data_valid    ( DownstreamStackBusLane[14][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane25_strm0_ready         ( DownstreamStackBusLane[14][25].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane25_strm0_cntl          ( DownstreamStackBusLane[14][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane25_strm0_data          ( DownstreamStackBusLane[14][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane25_strm0_data_valid    ( DownstreamStackBusLane[14][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane25_strm1_ready         ( DownstreamStackBusLane[14][25].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane25_strm1_cntl          ( DownstreamStackBusLane[14][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane25_strm1_data          ( DownstreamStackBusLane[14][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane25_strm1_data_valid    ( DownstreamStackBusLane[14][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane26_strm0_ready         ( DownstreamStackBusLane[14][26].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane26_strm0_cntl          ( DownstreamStackBusLane[14][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane26_strm0_data          ( DownstreamStackBusLane[14][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane26_strm0_data_valid    ( DownstreamStackBusLane[14][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane26_strm1_ready         ( DownstreamStackBusLane[14][26].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane26_strm1_cntl          ( DownstreamStackBusLane[14][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane26_strm1_data          ( DownstreamStackBusLane[14][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane26_strm1_data_valid    ( DownstreamStackBusLane[14][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane27_strm0_ready         ( DownstreamStackBusLane[14][27].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane27_strm0_cntl          ( DownstreamStackBusLane[14][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane27_strm0_data          ( DownstreamStackBusLane[14][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane27_strm0_data_valid    ( DownstreamStackBusLane[14][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane27_strm1_ready         ( DownstreamStackBusLane[14][27].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane27_strm1_cntl          ( DownstreamStackBusLane[14][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane27_strm1_data          ( DownstreamStackBusLane[14][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane27_strm1_data_valid    ( DownstreamStackBusLane[14][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane28_strm0_ready         ( DownstreamStackBusLane[14][28].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane28_strm0_cntl          ( DownstreamStackBusLane[14][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane28_strm0_data          ( DownstreamStackBusLane[14][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane28_strm0_data_valid    ( DownstreamStackBusLane[14][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane28_strm1_ready         ( DownstreamStackBusLane[14][28].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane28_strm1_cntl          ( DownstreamStackBusLane[14][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane28_strm1_data          ( DownstreamStackBusLane[14][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane28_strm1_data_valid    ( DownstreamStackBusLane[14][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane29_strm0_ready         ( DownstreamStackBusLane[14][29].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane29_strm0_cntl          ( DownstreamStackBusLane[14][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane29_strm0_data          ( DownstreamStackBusLane[14][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane29_strm0_data_valid    ( DownstreamStackBusLane[14][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane29_strm1_ready         ( DownstreamStackBusLane[14][29].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane29_strm1_cntl          ( DownstreamStackBusLane[14][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane29_strm1_data          ( DownstreamStackBusLane[14][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane29_strm1_data_valid    ( DownstreamStackBusLane[14][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane30_strm0_ready         ( DownstreamStackBusLane[14][30].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane30_strm0_cntl          ( DownstreamStackBusLane[14][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane30_strm0_data          ( DownstreamStackBusLane[14][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane30_strm0_data_valid    ( DownstreamStackBusLane[14][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane30_strm1_ready         ( DownstreamStackBusLane[14][30].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane30_strm1_cntl          ( DownstreamStackBusLane[14][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane30_strm1_data          ( DownstreamStackBusLane[14][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane30_strm1_data_valid    ( DownstreamStackBusLane[14][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 14, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane31_strm0_ready         ( DownstreamStackBusLane[14][31].pe__std__lane_strm0_ready              ),      
        .std__pe14__lane31_strm0_cntl          ( DownstreamStackBusLane[14][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe14__lane31_strm0_data          ( DownstreamStackBusLane[14][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe14__lane31_strm0_data_valid    ( DownstreamStackBusLane[14][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__std__lane31_strm1_ready         ( DownstreamStackBusLane[14][31].pe__std__lane_strm1_ready              ),      
        .std__pe14__lane31_strm1_cntl          ( DownstreamStackBusLane[14][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe14__lane31_strm1_data          ( DownstreamStackBusLane[14][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe14__lane31_strm1_data_valid    ( DownstreamStackBusLane[14][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane0_strm0_ready         ( DownstreamStackBusLane[15][0].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane0_strm0_cntl          ( DownstreamStackBusLane[15][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane0_strm0_data          ( DownstreamStackBusLane[15][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane0_strm0_data_valid    ( DownstreamStackBusLane[15][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane0_strm1_ready         ( DownstreamStackBusLane[15][0].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane0_strm1_cntl          ( DownstreamStackBusLane[15][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane0_strm1_data          ( DownstreamStackBusLane[15][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane0_strm1_data_valid    ( DownstreamStackBusLane[15][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane1_strm0_ready         ( DownstreamStackBusLane[15][1].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane1_strm0_cntl          ( DownstreamStackBusLane[15][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane1_strm0_data          ( DownstreamStackBusLane[15][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane1_strm0_data_valid    ( DownstreamStackBusLane[15][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane1_strm1_ready         ( DownstreamStackBusLane[15][1].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane1_strm1_cntl          ( DownstreamStackBusLane[15][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane1_strm1_data          ( DownstreamStackBusLane[15][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane1_strm1_data_valid    ( DownstreamStackBusLane[15][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane2_strm0_ready         ( DownstreamStackBusLane[15][2].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane2_strm0_cntl          ( DownstreamStackBusLane[15][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane2_strm0_data          ( DownstreamStackBusLane[15][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane2_strm0_data_valid    ( DownstreamStackBusLane[15][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane2_strm1_ready         ( DownstreamStackBusLane[15][2].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane2_strm1_cntl          ( DownstreamStackBusLane[15][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane2_strm1_data          ( DownstreamStackBusLane[15][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane2_strm1_data_valid    ( DownstreamStackBusLane[15][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane3_strm0_ready         ( DownstreamStackBusLane[15][3].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane3_strm0_cntl          ( DownstreamStackBusLane[15][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane3_strm0_data          ( DownstreamStackBusLane[15][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane3_strm0_data_valid    ( DownstreamStackBusLane[15][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane3_strm1_ready         ( DownstreamStackBusLane[15][3].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane3_strm1_cntl          ( DownstreamStackBusLane[15][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane3_strm1_data          ( DownstreamStackBusLane[15][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane3_strm1_data_valid    ( DownstreamStackBusLane[15][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane4_strm0_ready         ( DownstreamStackBusLane[15][4].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane4_strm0_cntl          ( DownstreamStackBusLane[15][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane4_strm0_data          ( DownstreamStackBusLane[15][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane4_strm0_data_valid    ( DownstreamStackBusLane[15][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane4_strm1_ready         ( DownstreamStackBusLane[15][4].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane4_strm1_cntl          ( DownstreamStackBusLane[15][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane4_strm1_data          ( DownstreamStackBusLane[15][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane4_strm1_data_valid    ( DownstreamStackBusLane[15][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane5_strm0_ready         ( DownstreamStackBusLane[15][5].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane5_strm0_cntl          ( DownstreamStackBusLane[15][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane5_strm0_data          ( DownstreamStackBusLane[15][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane5_strm0_data_valid    ( DownstreamStackBusLane[15][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane5_strm1_ready         ( DownstreamStackBusLane[15][5].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane5_strm1_cntl          ( DownstreamStackBusLane[15][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane5_strm1_data          ( DownstreamStackBusLane[15][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane5_strm1_data_valid    ( DownstreamStackBusLane[15][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane6_strm0_ready         ( DownstreamStackBusLane[15][6].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane6_strm0_cntl          ( DownstreamStackBusLane[15][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane6_strm0_data          ( DownstreamStackBusLane[15][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane6_strm0_data_valid    ( DownstreamStackBusLane[15][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane6_strm1_ready         ( DownstreamStackBusLane[15][6].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane6_strm1_cntl          ( DownstreamStackBusLane[15][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane6_strm1_data          ( DownstreamStackBusLane[15][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane6_strm1_data_valid    ( DownstreamStackBusLane[15][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane7_strm0_ready         ( DownstreamStackBusLane[15][7].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane7_strm0_cntl          ( DownstreamStackBusLane[15][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane7_strm0_data          ( DownstreamStackBusLane[15][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane7_strm0_data_valid    ( DownstreamStackBusLane[15][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane7_strm1_ready         ( DownstreamStackBusLane[15][7].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane7_strm1_cntl          ( DownstreamStackBusLane[15][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane7_strm1_data          ( DownstreamStackBusLane[15][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane7_strm1_data_valid    ( DownstreamStackBusLane[15][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane8_strm0_ready         ( DownstreamStackBusLane[15][8].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane8_strm0_cntl          ( DownstreamStackBusLane[15][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane8_strm0_data          ( DownstreamStackBusLane[15][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane8_strm0_data_valid    ( DownstreamStackBusLane[15][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane8_strm1_ready         ( DownstreamStackBusLane[15][8].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane8_strm1_cntl          ( DownstreamStackBusLane[15][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane8_strm1_data          ( DownstreamStackBusLane[15][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane8_strm1_data_valid    ( DownstreamStackBusLane[15][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane9_strm0_ready         ( DownstreamStackBusLane[15][9].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane9_strm0_cntl          ( DownstreamStackBusLane[15][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane9_strm0_data          ( DownstreamStackBusLane[15][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane9_strm0_data_valid    ( DownstreamStackBusLane[15][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane9_strm1_ready         ( DownstreamStackBusLane[15][9].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane9_strm1_cntl          ( DownstreamStackBusLane[15][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane9_strm1_data          ( DownstreamStackBusLane[15][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane9_strm1_data_valid    ( DownstreamStackBusLane[15][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane10_strm0_ready         ( DownstreamStackBusLane[15][10].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane10_strm0_cntl          ( DownstreamStackBusLane[15][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane10_strm0_data          ( DownstreamStackBusLane[15][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane10_strm0_data_valid    ( DownstreamStackBusLane[15][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane10_strm1_ready         ( DownstreamStackBusLane[15][10].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane10_strm1_cntl          ( DownstreamStackBusLane[15][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane10_strm1_data          ( DownstreamStackBusLane[15][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane10_strm1_data_valid    ( DownstreamStackBusLane[15][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane11_strm0_ready         ( DownstreamStackBusLane[15][11].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane11_strm0_cntl          ( DownstreamStackBusLane[15][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane11_strm0_data          ( DownstreamStackBusLane[15][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane11_strm0_data_valid    ( DownstreamStackBusLane[15][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane11_strm1_ready         ( DownstreamStackBusLane[15][11].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane11_strm1_cntl          ( DownstreamStackBusLane[15][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane11_strm1_data          ( DownstreamStackBusLane[15][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane11_strm1_data_valid    ( DownstreamStackBusLane[15][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane12_strm0_ready         ( DownstreamStackBusLane[15][12].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane12_strm0_cntl          ( DownstreamStackBusLane[15][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane12_strm0_data          ( DownstreamStackBusLane[15][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane12_strm0_data_valid    ( DownstreamStackBusLane[15][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane12_strm1_ready         ( DownstreamStackBusLane[15][12].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane12_strm1_cntl          ( DownstreamStackBusLane[15][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane12_strm1_data          ( DownstreamStackBusLane[15][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane12_strm1_data_valid    ( DownstreamStackBusLane[15][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane13_strm0_ready         ( DownstreamStackBusLane[15][13].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane13_strm0_cntl          ( DownstreamStackBusLane[15][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane13_strm0_data          ( DownstreamStackBusLane[15][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane13_strm0_data_valid    ( DownstreamStackBusLane[15][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane13_strm1_ready         ( DownstreamStackBusLane[15][13].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane13_strm1_cntl          ( DownstreamStackBusLane[15][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane13_strm1_data          ( DownstreamStackBusLane[15][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane13_strm1_data_valid    ( DownstreamStackBusLane[15][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane14_strm0_ready         ( DownstreamStackBusLane[15][14].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane14_strm0_cntl          ( DownstreamStackBusLane[15][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane14_strm0_data          ( DownstreamStackBusLane[15][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane14_strm0_data_valid    ( DownstreamStackBusLane[15][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane14_strm1_ready         ( DownstreamStackBusLane[15][14].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane14_strm1_cntl          ( DownstreamStackBusLane[15][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane14_strm1_data          ( DownstreamStackBusLane[15][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane14_strm1_data_valid    ( DownstreamStackBusLane[15][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane15_strm0_ready         ( DownstreamStackBusLane[15][15].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane15_strm0_cntl          ( DownstreamStackBusLane[15][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane15_strm0_data          ( DownstreamStackBusLane[15][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane15_strm0_data_valid    ( DownstreamStackBusLane[15][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane15_strm1_ready         ( DownstreamStackBusLane[15][15].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane15_strm1_cntl          ( DownstreamStackBusLane[15][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane15_strm1_data          ( DownstreamStackBusLane[15][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane15_strm1_data_valid    ( DownstreamStackBusLane[15][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane16_strm0_ready         ( DownstreamStackBusLane[15][16].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane16_strm0_cntl          ( DownstreamStackBusLane[15][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane16_strm0_data          ( DownstreamStackBusLane[15][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane16_strm0_data_valid    ( DownstreamStackBusLane[15][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane16_strm1_ready         ( DownstreamStackBusLane[15][16].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane16_strm1_cntl          ( DownstreamStackBusLane[15][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane16_strm1_data          ( DownstreamStackBusLane[15][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane16_strm1_data_valid    ( DownstreamStackBusLane[15][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane17_strm0_ready         ( DownstreamStackBusLane[15][17].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane17_strm0_cntl          ( DownstreamStackBusLane[15][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane17_strm0_data          ( DownstreamStackBusLane[15][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane17_strm0_data_valid    ( DownstreamStackBusLane[15][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane17_strm1_ready         ( DownstreamStackBusLane[15][17].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane17_strm1_cntl          ( DownstreamStackBusLane[15][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane17_strm1_data          ( DownstreamStackBusLane[15][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane17_strm1_data_valid    ( DownstreamStackBusLane[15][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane18_strm0_ready         ( DownstreamStackBusLane[15][18].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane18_strm0_cntl          ( DownstreamStackBusLane[15][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane18_strm0_data          ( DownstreamStackBusLane[15][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane18_strm0_data_valid    ( DownstreamStackBusLane[15][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane18_strm1_ready         ( DownstreamStackBusLane[15][18].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane18_strm1_cntl          ( DownstreamStackBusLane[15][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane18_strm1_data          ( DownstreamStackBusLane[15][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane18_strm1_data_valid    ( DownstreamStackBusLane[15][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane19_strm0_ready         ( DownstreamStackBusLane[15][19].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane19_strm0_cntl          ( DownstreamStackBusLane[15][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane19_strm0_data          ( DownstreamStackBusLane[15][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane19_strm0_data_valid    ( DownstreamStackBusLane[15][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane19_strm1_ready         ( DownstreamStackBusLane[15][19].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane19_strm1_cntl          ( DownstreamStackBusLane[15][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane19_strm1_data          ( DownstreamStackBusLane[15][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane19_strm1_data_valid    ( DownstreamStackBusLane[15][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane20_strm0_ready         ( DownstreamStackBusLane[15][20].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane20_strm0_cntl          ( DownstreamStackBusLane[15][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane20_strm0_data          ( DownstreamStackBusLane[15][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane20_strm0_data_valid    ( DownstreamStackBusLane[15][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane20_strm1_ready         ( DownstreamStackBusLane[15][20].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane20_strm1_cntl          ( DownstreamStackBusLane[15][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane20_strm1_data          ( DownstreamStackBusLane[15][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane20_strm1_data_valid    ( DownstreamStackBusLane[15][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane21_strm0_ready         ( DownstreamStackBusLane[15][21].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane21_strm0_cntl          ( DownstreamStackBusLane[15][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane21_strm0_data          ( DownstreamStackBusLane[15][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane21_strm0_data_valid    ( DownstreamStackBusLane[15][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane21_strm1_ready         ( DownstreamStackBusLane[15][21].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane21_strm1_cntl          ( DownstreamStackBusLane[15][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane21_strm1_data          ( DownstreamStackBusLane[15][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane21_strm1_data_valid    ( DownstreamStackBusLane[15][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane22_strm0_ready         ( DownstreamStackBusLane[15][22].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane22_strm0_cntl          ( DownstreamStackBusLane[15][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane22_strm0_data          ( DownstreamStackBusLane[15][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane22_strm0_data_valid    ( DownstreamStackBusLane[15][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane22_strm1_ready         ( DownstreamStackBusLane[15][22].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane22_strm1_cntl          ( DownstreamStackBusLane[15][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane22_strm1_data          ( DownstreamStackBusLane[15][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane22_strm1_data_valid    ( DownstreamStackBusLane[15][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane23_strm0_ready         ( DownstreamStackBusLane[15][23].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane23_strm0_cntl          ( DownstreamStackBusLane[15][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane23_strm0_data          ( DownstreamStackBusLane[15][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane23_strm0_data_valid    ( DownstreamStackBusLane[15][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane23_strm1_ready         ( DownstreamStackBusLane[15][23].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane23_strm1_cntl          ( DownstreamStackBusLane[15][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane23_strm1_data          ( DownstreamStackBusLane[15][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane23_strm1_data_valid    ( DownstreamStackBusLane[15][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane24_strm0_ready         ( DownstreamStackBusLane[15][24].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane24_strm0_cntl          ( DownstreamStackBusLane[15][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane24_strm0_data          ( DownstreamStackBusLane[15][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane24_strm0_data_valid    ( DownstreamStackBusLane[15][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane24_strm1_ready         ( DownstreamStackBusLane[15][24].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane24_strm1_cntl          ( DownstreamStackBusLane[15][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane24_strm1_data          ( DownstreamStackBusLane[15][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane24_strm1_data_valid    ( DownstreamStackBusLane[15][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane25_strm0_ready         ( DownstreamStackBusLane[15][25].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane25_strm0_cntl          ( DownstreamStackBusLane[15][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane25_strm0_data          ( DownstreamStackBusLane[15][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane25_strm0_data_valid    ( DownstreamStackBusLane[15][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane25_strm1_ready         ( DownstreamStackBusLane[15][25].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane25_strm1_cntl          ( DownstreamStackBusLane[15][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane25_strm1_data          ( DownstreamStackBusLane[15][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane25_strm1_data_valid    ( DownstreamStackBusLane[15][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane26_strm0_ready         ( DownstreamStackBusLane[15][26].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane26_strm0_cntl          ( DownstreamStackBusLane[15][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane26_strm0_data          ( DownstreamStackBusLane[15][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane26_strm0_data_valid    ( DownstreamStackBusLane[15][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane26_strm1_ready         ( DownstreamStackBusLane[15][26].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane26_strm1_cntl          ( DownstreamStackBusLane[15][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane26_strm1_data          ( DownstreamStackBusLane[15][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane26_strm1_data_valid    ( DownstreamStackBusLane[15][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane27_strm0_ready         ( DownstreamStackBusLane[15][27].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane27_strm0_cntl          ( DownstreamStackBusLane[15][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane27_strm0_data          ( DownstreamStackBusLane[15][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane27_strm0_data_valid    ( DownstreamStackBusLane[15][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane27_strm1_ready         ( DownstreamStackBusLane[15][27].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane27_strm1_cntl          ( DownstreamStackBusLane[15][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane27_strm1_data          ( DownstreamStackBusLane[15][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane27_strm1_data_valid    ( DownstreamStackBusLane[15][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane28_strm0_ready         ( DownstreamStackBusLane[15][28].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane28_strm0_cntl          ( DownstreamStackBusLane[15][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane28_strm0_data          ( DownstreamStackBusLane[15][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane28_strm0_data_valid    ( DownstreamStackBusLane[15][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane28_strm1_ready         ( DownstreamStackBusLane[15][28].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane28_strm1_cntl          ( DownstreamStackBusLane[15][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane28_strm1_data          ( DownstreamStackBusLane[15][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane28_strm1_data_valid    ( DownstreamStackBusLane[15][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane29_strm0_ready         ( DownstreamStackBusLane[15][29].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane29_strm0_cntl          ( DownstreamStackBusLane[15][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane29_strm0_data          ( DownstreamStackBusLane[15][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane29_strm0_data_valid    ( DownstreamStackBusLane[15][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane29_strm1_ready         ( DownstreamStackBusLane[15][29].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane29_strm1_cntl          ( DownstreamStackBusLane[15][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane29_strm1_data          ( DownstreamStackBusLane[15][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane29_strm1_data_valid    ( DownstreamStackBusLane[15][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane30_strm0_ready         ( DownstreamStackBusLane[15][30].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane30_strm0_cntl          ( DownstreamStackBusLane[15][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane30_strm0_data          ( DownstreamStackBusLane[15][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane30_strm0_data_valid    ( DownstreamStackBusLane[15][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane30_strm1_ready         ( DownstreamStackBusLane[15][30].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane30_strm1_cntl          ( DownstreamStackBusLane[15][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane30_strm1_data          ( DownstreamStackBusLane[15][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane30_strm1_data_valid    ( DownstreamStackBusLane[15][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 15, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane31_strm0_ready         ( DownstreamStackBusLane[15][31].pe__std__lane_strm0_ready              ),      
        .std__pe15__lane31_strm0_cntl          ( DownstreamStackBusLane[15][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe15__lane31_strm0_data          ( DownstreamStackBusLane[15][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe15__lane31_strm0_data_valid    ( DownstreamStackBusLane[15][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__std__lane31_strm1_ready         ( DownstreamStackBusLane[15][31].pe__std__lane_strm1_ready              ),      
        .std__pe15__lane31_strm1_cntl          ( DownstreamStackBusLane[15][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe15__lane31_strm1_data          ( DownstreamStackBusLane[15][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe15__lane31_strm1_data_valid    ( DownstreamStackBusLane[15][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane0_strm0_ready         ( DownstreamStackBusLane[16][0].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane0_strm0_cntl          ( DownstreamStackBusLane[16][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane0_strm0_data          ( DownstreamStackBusLane[16][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane0_strm0_data_valid    ( DownstreamStackBusLane[16][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane0_strm1_ready         ( DownstreamStackBusLane[16][0].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane0_strm1_cntl          ( DownstreamStackBusLane[16][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane0_strm1_data          ( DownstreamStackBusLane[16][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane0_strm1_data_valid    ( DownstreamStackBusLane[16][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane1_strm0_ready         ( DownstreamStackBusLane[16][1].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane1_strm0_cntl          ( DownstreamStackBusLane[16][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane1_strm0_data          ( DownstreamStackBusLane[16][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane1_strm0_data_valid    ( DownstreamStackBusLane[16][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane1_strm1_ready         ( DownstreamStackBusLane[16][1].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane1_strm1_cntl          ( DownstreamStackBusLane[16][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane1_strm1_data          ( DownstreamStackBusLane[16][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane1_strm1_data_valid    ( DownstreamStackBusLane[16][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane2_strm0_ready         ( DownstreamStackBusLane[16][2].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane2_strm0_cntl          ( DownstreamStackBusLane[16][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane2_strm0_data          ( DownstreamStackBusLane[16][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane2_strm0_data_valid    ( DownstreamStackBusLane[16][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane2_strm1_ready         ( DownstreamStackBusLane[16][2].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane2_strm1_cntl          ( DownstreamStackBusLane[16][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane2_strm1_data          ( DownstreamStackBusLane[16][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane2_strm1_data_valid    ( DownstreamStackBusLane[16][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane3_strm0_ready         ( DownstreamStackBusLane[16][3].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane3_strm0_cntl          ( DownstreamStackBusLane[16][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane3_strm0_data          ( DownstreamStackBusLane[16][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane3_strm0_data_valid    ( DownstreamStackBusLane[16][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane3_strm1_ready         ( DownstreamStackBusLane[16][3].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane3_strm1_cntl          ( DownstreamStackBusLane[16][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane3_strm1_data          ( DownstreamStackBusLane[16][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane3_strm1_data_valid    ( DownstreamStackBusLane[16][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane4_strm0_ready         ( DownstreamStackBusLane[16][4].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane4_strm0_cntl          ( DownstreamStackBusLane[16][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane4_strm0_data          ( DownstreamStackBusLane[16][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane4_strm0_data_valid    ( DownstreamStackBusLane[16][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane4_strm1_ready         ( DownstreamStackBusLane[16][4].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane4_strm1_cntl          ( DownstreamStackBusLane[16][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane4_strm1_data          ( DownstreamStackBusLane[16][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane4_strm1_data_valid    ( DownstreamStackBusLane[16][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane5_strm0_ready         ( DownstreamStackBusLane[16][5].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane5_strm0_cntl          ( DownstreamStackBusLane[16][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane5_strm0_data          ( DownstreamStackBusLane[16][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane5_strm0_data_valid    ( DownstreamStackBusLane[16][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane5_strm1_ready         ( DownstreamStackBusLane[16][5].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane5_strm1_cntl          ( DownstreamStackBusLane[16][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane5_strm1_data          ( DownstreamStackBusLane[16][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane5_strm1_data_valid    ( DownstreamStackBusLane[16][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane6_strm0_ready         ( DownstreamStackBusLane[16][6].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane6_strm0_cntl          ( DownstreamStackBusLane[16][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane6_strm0_data          ( DownstreamStackBusLane[16][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane6_strm0_data_valid    ( DownstreamStackBusLane[16][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane6_strm1_ready         ( DownstreamStackBusLane[16][6].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane6_strm1_cntl          ( DownstreamStackBusLane[16][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane6_strm1_data          ( DownstreamStackBusLane[16][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane6_strm1_data_valid    ( DownstreamStackBusLane[16][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane7_strm0_ready         ( DownstreamStackBusLane[16][7].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane7_strm0_cntl          ( DownstreamStackBusLane[16][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane7_strm0_data          ( DownstreamStackBusLane[16][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane7_strm0_data_valid    ( DownstreamStackBusLane[16][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane7_strm1_ready         ( DownstreamStackBusLane[16][7].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane7_strm1_cntl          ( DownstreamStackBusLane[16][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane7_strm1_data          ( DownstreamStackBusLane[16][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane7_strm1_data_valid    ( DownstreamStackBusLane[16][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane8_strm0_ready         ( DownstreamStackBusLane[16][8].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane8_strm0_cntl          ( DownstreamStackBusLane[16][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane8_strm0_data          ( DownstreamStackBusLane[16][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane8_strm0_data_valid    ( DownstreamStackBusLane[16][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane8_strm1_ready         ( DownstreamStackBusLane[16][8].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane8_strm1_cntl          ( DownstreamStackBusLane[16][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane8_strm1_data          ( DownstreamStackBusLane[16][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane8_strm1_data_valid    ( DownstreamStackBusLane[16][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane9_strm0_ready         ( DownstreamStackBusLane[16][9].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane9_strm0_cntl          ( DownstreamStackBusLane[16][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane9_strm0_data          ( DownstreamStackBusLane[16][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane9_strm0_data_valid    ( DownstreamStackBusLane[16][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane9_strm1_ready         ( DownstreamStackBusLane[16][9].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane9_strm1_cntl          ( DownstreamStackBusLane[16][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane9_strm1_data          ( DownstreamStackBusLane[16][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane9_strm1_data_valid    ( DownstreamStackBusLane[16][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane10_strm0_ready         ( DownstreamStackBusLane[16][10].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane10_strm0_cntl          ( DownstreamStackBusLane[16][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane10_strm0_data          ( DownstreamStackBusLane[16][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane10_strm0_data_valid    ( DownstreamStackBusLane[16][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane10_strm1_ready         ( DownstreamStackBusLane[16][10].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane10_strm1_cntl          ( DownstreamStackBusLane[16][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane10_strm1_data          ( DownstreamStackBusLane[16][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane10_strm1_data_valid    ( DownstreamStackBusLane[16][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane11_strm0_ready         ( DownstreamStackBusLane[16][11].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane11_strm0_cntl          ( DownstreamStackBusLane[16][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane11_strm0_data          ( DownstreamStackBusLane[16][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane11_strm0_data_valid    ( DownstreamStackBusLane[16][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane11_strm1_ready         ( DownstreamStackBusLane[16][11].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane11_strm1_cntl          ( DownstreamStackBusLane[16][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane11_strm1_data          ( DownstreamStackBusLane[16][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane11_strm1_data_valid    ( DownstreamStackBusLane[16][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane12_strm0_ready         ( DownstreamStackBusLane[16][12].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane12_strm0_cntl          ( DownstreamStackBusLane[16][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane12_strm0_data          ( DownstreamStackBusLane[16][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane12_strm0_data_valid    ( DownstreamStackBusLane[16][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane12_strm1_ready         ( DownstreamStackBusLane[16][12].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane12_strm1_cntl          ( DownstreamStackBusLane[16][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane12_strm1_data          ( DownstreamStackBusLane[16][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane12_strm1_data_valid    ( DownstreamStackBusLane[16][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane13_strm0_ready         ( DownstreamStackBusLane[16][13].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane13_strm0_cntl          ( DownstreamStackBusLane[16][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane13_strm0_data          ( DownstreamStackBusLane[16][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane13_strm0_data_valid    ( DownstreamStackBusLane[16][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane13_strm1_ready         ( DownstreamStackBusLane[16][13].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane13_strm1_cntl          ( DownstreamStackBusLane[16][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane13_strm1_data          ( DownstreamStackBusLane[16][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane13_strm1_data_valid    ( DownstreamStackBusLane[16][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane14_strm0_ready         ( DownstreamStackBusLane[16][14].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane14_strm0_cntl          ( DownstreamStackBusLane[16][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane14_strm0_data          ( DownstreamStackBusLane[16][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane14_strm0_data_valid    ( DownstreamStackBusLane[16][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane14_strm1_ready         ( DownstreamStackBusLane[16][14].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane14_strm1_cntl          ( DownstreamStackBusLane[16][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane14_strm1_data          ( DownstreamStackBusLane[16][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane14_strm1_data_valid    ( DownstreamStackBusLane[16][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane15_strm0_ready         ( DownstreamStackBusLane[16][15].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane15_strm0_cntl          ( DownstreamStackBusLane[16][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane15_strm0_data          ( DownstreamStackBusLane[16][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane15_strm0_data_valid    ( DownstreamStackBusLane[16][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane15_strm1_ready         ( DownstreamStackBusLane[16][15].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane15_strm1_cntl          ( DownstreamStackBusLane[16][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane15_strm1_data          ( DownstreamStackBusLane[16][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane15_strm1_data_valid    ( DownstreamStackBusLane[16][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane16_strm0_ready         ( DownstreamStackBusLane[16][16].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane16_strm0_cntl          ( DownstreamStackBusLane[16][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane16_strm0_data          ( DownstreamStackBusLane[16][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane16_strm0_data_valid    ( DownstreamStackBusLane[16][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane16_strm1_ready         ( DownstreamStackBusLane[16][16].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane16_strm1_cntl          ( DownstreamStackBusLane[16][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane16_strm1_data          ( DownstreamStackBusLane[16][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane16_strm1_data_valid    ( DownstreamStackBusLane[16][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane17_strm0_ready         ( DownstreamStackBusLane[16][17].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane17_strm0_cntl          ( DownstreamStackBusLane[16][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane17_strm0_data          ( DownstreamStackBusLane[16][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane17_strm0_data_valid    ( DownstreamStackBusLane[16][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane17_strm1_ready         ( DownstreamStackBusLane[16][17].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane17_strm1_cntl          ( DownstreamStackBusLane[16][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane17_strm1_data          ( DownstreamStackBusLane[16][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane17_strm1_data_valid    ( DownstreamStackBusLane[16][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane18_strm0_ready         ( DownstreamStackBusLane[16][18].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane18_strm0_cntl          ( DownstreamStackBusLane[16][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane18_strm0_data          ( DownstreamStackBusLane[16][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane18_strm0_data_valid    ( DownstreamStackBusLane[16][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane18_strm1_ready         ( DownstreamStackBusLane[16][18].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane18_strm1_cntl          ( DownstreamStackBusLane[16][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane18_strm1_data          ( DownstreamStackBusLane[16][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane18_strm1_data_valid    ( DownstreamStackBusLane[16][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane19_strm0_ready         ( DownstreamStackBusLane[16][19].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane19_strm0_cntl          ( DownstreamStackBusLane[16][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane19_strm0_data          ( DownstreamStackBusLane[16][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane19_strm0_data_valid    ( DownstreamStackBusLane[16][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane19_strm1_ready         ( DownstreamStackBusLane[16][19].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane19_strm1_cntl          ( DownstreamStackBusLane[16][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane19_strm1_data          ( DownstreamStackBusLane[16][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane19_strm1_data_valid    ( DownstreamStackBusLane[16][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane20_strm0_ready         ( DownstreamStackBusLane[16][20].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane20_strm0_cntl          ( DownstreamStackBusLane[16][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane20_strm0_data          ( DownstreamStackBusLane[16][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane20_strm0_data_valid    ( DownstreamStackBusLane[16][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane20_strm1_ready         ( DownstreamStackBusLane[16][20].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane20_strm1_cntl          ( DownstreamStackBusLane[16][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane20_strm1_data          ( DownstreamStackBusLane[16][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane20_strm1_data_valid    ( DownstreamStackBusLane[16][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane21_strm0_ready         ( DownstreamStackBusLane[16][21].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane21_strm0_cntl          ( DownstreamStackBusLane[16][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane21_strm0_data          ( DownstreamStackBusLane[16][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane21_strm0_data_valid    ( DownstreamStackBusLane[16][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane21_strm1_ready         ( DownstreamStackBusLane[16][21].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane21_strm1_cntl          ( DownstreamStackBusLane[16][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane21_strm1_data          ( DownstreamStackBusLane[16][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane21_strm1_data_valid    ( DownstreamStackBusLane[16][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane22_strm0_ready         ( DownstreamStackBusLane[16][22].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane22_strm0_cntl          ( DownstreamStackBusLane[16][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane22_strm0_data          ( DownstreamStackBusLane[16][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane22_strm0_data_valid    ( DownstreamStackBusLane[16][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane22_strm1_ready         ( DownstreamStackBusLane[16][22].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane22_strm1_cntl          ( DownstreamStackBusLane[16][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane22_strm1_data          ( DownstreamStackBusLane[16][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane22_strm1_data_valid    ( DownstreamStackBusLane[16][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane23_strm0_ready         ( DownstreamStackBusLane[16][23].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane23_strm0_cntl          ( DownstreamStackBusLane[16][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane23_strm0_data          ( DownstreamStackBusLane[16][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane23_strm0_data_valid    ( DownstreamStackBusLane[16][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane23_strm1_ready         ( DownstreamStackBusLane[16][23].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane23_strm1_cntl          ( DownstreamStackBusLane[16][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane23_strm1_data          ( DownstreamStackBusLane[16][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane23_strm1_data_valid    ( DownstreamStackBusLane[16][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane24_strm0_ready         ( DownstreamStackBusLane[16][24].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane24_strm0_cntl          ( DownstreamStackBusLane[16][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane24_strm0_data          ( DownstreamStackBusLane[16][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane24_strm0_data_valid    ( DownstreamStackBusLane[16][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane24_strm1_ready         ( DownstreamStackBusLane[16][24].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane24_strm1_cntl          ( DownstreamStackBusLane[16][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane24_strm1_data          ( DownstreamStackBusLane[16][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane24_strm1_data_valid    ( DownstreamStackBusLane[16][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane25_strm0_ready         ( DownstreamStackBusLane[16][25].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane25_strm0_cntl          ( DownstreamStackBusLane[16][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane25_strm0_data          ( DownstreamStackBusLane[16][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane25_strm0_data_valid    ( DownstreamStackBusLane[16][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane25_strm1_ready         ( DownstreamStackBusLane[16][25].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane25_strm1_cntl          ( DownstreamStackBusLane[16][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane25_strm1_data          ( DownstreamStackBusLane[16][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane25_strm1_data_valid    ( DownstreamStackBusLane[16][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane26_strm0_ready         ( DownstreamStackBusLane[16][26].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane26_strm0_cntl          ( DownstreamStackBusLane[16][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane26_strm0_data          ( DownstreamStackBusLane[16][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane26_strm0_data_valid    ( DownstreamStackBusLane[16][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane26_strm1_ready         ( DownstreamStackBusLane[16][26].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane26_strm1_cntl          ( DownstreamStackBusLane[16][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane26_strm1_data          ( DownstreamStackBusLane[16][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane26_strm1_data_valid    ( DownstreamStackBusLane[16][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane27_strm0_ready         ( DownstreamStackBusLane[16][27].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane27_strm0_cntl          ( DownstreamStackBusLane[16][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane27_strm0_data          ( DownstreamStackBusLane[16][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane27_strm0_data_valid    ( DownstreamStackBusLane[16][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane27_strm1_ready         ( DownstreamStackBusLane[16][27].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane27_strm1_cntl          ( DownstreamStackBusLane[16][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane27_strm1_data          ( DownstreamStackBusLane[16][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane27_strm1_data_valid    ( DownstreamStackBusLane[16][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane28_strm0_ready         ( DownstreamStackBusLane[16][28].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane28_strm0_cntl          ( DownstreamStackBusLane[16][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane28_strm0_data          ( DownstreamStackBusLane[16][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane28_strm0_data_valid    ( DownstreamStackBusLane[16][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane28_strm1_ready         ( DownstreamStackBusLane[16][28].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane28_strm1_cntl          ( DownstreamStackBusLane[16][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane28_strm1_data          ( DownstreamStackBusLane[16][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane28_strm1_data_valid    ( DownstreamStackBusLane[16][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane29_strm0_ready         ( DownstreamStackBusLane[16][29].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane29_strm0_cntl          ( DownstreamStackBusLane[16][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane29_strm0_data          ( DownstreamStackBusLane[16][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane29_strm0_data_valid    ( DownstreamStackBusLane[16][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane29_strm1_ready         ( DownstreamStackBusLane[16][29].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane29_strm1_cntl          ( DownstreamStackBusLane[16][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane29_strm1_data          ( DownstreamStackBusLane[16][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane29_strm1_data_valid    ( DownstreamStackBusLane[16][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane30_strm0_ready         ( DownstreamStackBusLane[16][30].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane30_strm0_cntl          ( DownstreamStackBusLane[16][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane30_strm0_data          ( DownstreamStackBusLane[16][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane30_strm0_data_valid    ( DownstreamStackBusLane[16][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane30_strm1_ready         ( DownstreamStackBusLane[16][30].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane30_strm1_cntl          ( DownstreamStackBusLane[16][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane30_strm1_data          ( DownstreamStackBusLane[16][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane30_strm1_data_valid    ( DownstreamStackBusLane[16][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 16, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane31_strm0_ready         ( DownstreamStackBusLane[16][31].pe__std__lane_strm0_ready              ),      
        .std__pe16__lane31_strm0_cntl          ( DownstreamStackBusLane[16][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe16__lane31_strm0_data          ( DownstreamStackBusLane[16][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe16__lane31_strm0_data_valid    ( DownstreamStackBusLane[16][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__std__lane31_strm1_ready         ( DownstreamStackBusLane[16][31].pe__std__lane_strm1_ready              ),      
        .std__pe16__lane31_strm1_cntl          ( DownstreamStackBusLane[16][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe16__lane31_strm1_data          ( DownstreamStackBusLane[16][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe16__lane31_strm1_data_valid    ( DownstreamStackBusLane[16][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane0_strm0_ready         ( DownstreamStackBusLane[17][0].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane0_strm0_cntl          ( DownstreamStackBusLane[17][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane0_strm0_data          ( DownstreamStackBusLane[17][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane0_strm0_data_valid    ( DownstreamStackBusLane[17][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane0_strm1_ready         ( DownstreamStackBusLane[17][0].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane0_strm1_cntl          ( DownstreamStackBusLane[17][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane0_strm1_data          ( DownstreamStackBusLane[17][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane0_strm1_data_valid    ( DownstreamStackBusLane[17][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane1_strm0_ready         ( DownstreamStackBusLane[17][1].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane1_strm0_cntl          ( DownstreamStackBusLane[17][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane1_strm0_data          ( DownstreamStackBusLane[17][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane1_strm0_data_valid    ( DownstreamStackBusLane[17][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane1_strm1_ready         ( DownstreamStackBusLane[17][1].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane1_strm1_cntl          ( DownstreamStackBusLane[17][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane1_strm1_data          ( DownstreamStackBusLane[17][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane1_strm1_data_valid    ( DownstreamStackBusLane[17][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane2_strm0_ready         ( DownstreamStackBusLane[17][2].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane2_strm0_cntl          ( DownstreamStackBusLane[17][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane2_strm0_data          ( DownstreamStackBusLane[17][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane2_strm0_data_valid    ( DownstreamStackBusLane[17][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane2_strm1_ready         ( DownstreamStackBusLane[17][2].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane2_strm1_cntl          ( DownstreamStackBusLane[17][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane2_strm1_data          ( DownstreamStackBusLane[17][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane2_strm1_data_valid    ( DownstreamStackBusLane[17][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane3_strm0_ready         ( DownstreamStackBusLane[17][3].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane3_strm0_cntl          ( DownstreamStackBusLane[17][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane3_strm0_data          ( DownstreamStackBusLane[17][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane3_strm0_data_valid    ( DownstreamStackBusLane[17][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane3_strm1_ready         ( DownstreamStackBusLane[17][3].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane3_strm1_cntl          ( DownstreamStackBusLane[17][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane3_strm1_data          ( DownstreamStackBusLane[17][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane3_strm1_data_valid    ( DownstreamStackBusLane[17][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane4_strm0_ready         ( DownstreamStackBusLane[17][4].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane4_strm0_cntl          ( DownstreamStackBusLane[17][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane4_strm0_data          ( DownstreamStackBusLane[17][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane4_strm0_data_valid    ( DownstreamStackBusLane[17][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane4_strm1_ready         ( DownstreamStackBusLane[17][4].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane4_strm1_cntl          ( DownstreamStackBusLane[17][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane4_strm1_data          ( DownstreamStackBusLane[17][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane4_strm1_data_valid    ( DownstreamStackBusLane[17][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane5_strm0_ready         ( DownstreamStackBusLane[17][5].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane5_strm0_cntl          ( DownstreamStackBusLane[17][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane5_strm0_data          ( DownstreamStackBusLane[17][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane5_strm0_data_valid    ( DownstreamStackBusLane[17][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane5_strm1_ready         ( DownstreamStackBusLane[17][5].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane5_strm1_cntl          ( DownstreamStackBusLane[17][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane5_strm1_data          ( DownstreamStackBusLane[17][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane5_strm1_data_valid    ( DownstreamStackBusLane[17][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane6_strm0_ready         ( DownstreamStackBusLane[17][6].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane6_strm0_cntl          ( DownstreamStackBusLane[17][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane6_strm0_data          ( DownstreamStackBusLane[17][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane6_strm0_data_valid    ( DownstreamStackBusLane[17][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane6_strm1_ready         ( DownstreamStackBusLane[17][6].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane6_strm1_cntl          ( DownstreamStackBusLane[17][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane6_strm1_data          ( DownstreamStackBusLane[17][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane6_strm1_data_valid    ( DownstreamStackBusLane[17][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane7_strm0_ready         ( DownstreamStackBusLane[17][7].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane7_strm0_cntl          ( DownstreamStackBusLane[17][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane7_strm0_data          ( DownstreamStackBusLane[17][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane7_strm0_data_valid    ( DownstreamStackBusLane[17][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane7_strm1_ready         ( DownstreamStackBusLane[17][7].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane7_strm1_cntl          ( DownstreamStackBusLane[17][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane7_strm1_data          ( DownstreamStackBusLane[17][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane7_strm1_data_valid    ( DownstreamStackBusLane[17][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane8_strm0_ready         ( DownstreamStackBusLane[17][8].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane8_strm0_cntl          ( DownstreamStackBusLane[17][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane8_strm0_data          ( DownstreamStackBusLane[17][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane8_strm0_data_valid    ( DownstreamStackBusLane[17][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane8_strm1_ready         ( DownstreamStackBusLane[17][8].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane8_strm1_cntl          ( DownstreamStackBusLane[17][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane8_strm1_data          ( DownstreamStackBusLane[17][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane8_strm1_data_valid    ( DownstreamStackBusLane[17][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane9_strm0_ready         ( DownstreamStackBusLane[17][9].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane9_strm0_cntl          ( DownstreamStackBusLane[17][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane9_strm0_data          ( DownstreamStackBusLane[17][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane9_strm0_data_valid    ( DownstreamStackBusLane[17][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane9_strm1_ready         ( DownstreamStackBusLane[17][9].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane9_strm1_cntl          ( DownstreamStackBusLane[17][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane9_strm1_data          ( DownstreamStackBusLane[17][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane9_strm1_data_valid    ( DownstreamStackBusLane[17][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane10_strm0_ready         ( DownstreamStackBusLane[17][10].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane10_strm0_cntl          ( DownstreamStackBusLane[17][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane10_strm0_data          ( DownstreamStackBusLane[17][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane10_strm0_data_valid    ( DownstreamStackBusLane[17][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane10_strm1_ready         ( DownstreamStackBusLane[17][10].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane10_strm1_cntl          ( DownstreamStackBusLane[17][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane10_strm1_data          ( DownstreamStackBusLane[17][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane10_strm1_data_valid    ( DownstreamStackBusLane[17][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane11_strm0_ready         ( DownstreamStackBusLane[17][11].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane11_strm0_cntl          ( DownstreamStackBusLane[17][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane11_strm0_data          ( DownstreamStackBusLane[17][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane11_strm0_data_valid    ( DownstreamStackBusLane[17][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane11_strm1_ready         ( DownstreamStackBusLane[17][11].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane11_strm1_cntl          ( DownstreamStackBusLane[17][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane11_strm1_data          ( DownstreamStackBusLane[17][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane11_strm1_data_valid    ( DownstreamStackBusLane[17][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane12_strm0_ready         ( DownstreamStackBusLane[17][12].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane12_strm0_cntl          ( DownstreamStackBusLane[17][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane12_strm0_data          ( DownstreamStackBusLane[17][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane12_strm0_data_valid    ( DownstreamStackBusLane[17][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane12_strm1_ready         ( DownstreamStackBusLane[17][12].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane12_strm1_cntl          ( DownstreamStackBusLane[17][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane12_strm1_data          ( DownstreamStackBusLane[17][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane12_strm1_data_valid    ( DownstreamStackBusLane[17][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane13_strm0_ready         ( DownstreamStackBusLane[17][13].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane13_strm0_cntl          ( DownstreamStackBusLane[17][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane13_strm0_data          ( DownstreamStackBusLane[17][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane13_strm0_data_valid    ( DownstreamStackBusLane[17][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane13_strm1_ready         ( DownstreamStackBusLane[17][13].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane13_strm1_cntl          ( DownstreamStackBusLane[17][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane13_strm1_data          ( DownstreamStackBusLane[17][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane13_strm1_data_valid    ( DownstreamStackBusLane[17][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane14_strm0_ready         ( DownstreamStackBusLane[17][14].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane14_strm0_cntl          ( DownstreamStackBusLane[17][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane14_strm0_data          ( DownstreamStackBusLane[17][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane14_strm0_data_valid    ( DownstreamStackBusLane[17][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane14_strm1_ready         ( DownstreamStackBusLane[17][14].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane14_strm1_cntl          ( DownstreamStackBusLane[17][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane14_strm1_data          ( DownstreamStackBusLane[17][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane14_strm1_data_valid    ( DownstreamStackBusLane[17][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane15_strm0_ready         ( DownstreamStackBusLane[17][15].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane15_strm0_cntl          ( DownstreamStackBusLane[17][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane15_strm0_data          ( DownstreamStackBusLane[17][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane15_strm0_data_valid    ( DownstreamStackBusLane[17][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane15_strm1_ready         ( DownstreamStackBusLane[17][15].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane15_strm1_cntl          ( DownstreamStackBusLane[17][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane15_strm1_data          ( DownstreamStackBusLane[17][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane15_strm1_data_valid    ( DownstreamStackBusLane[17][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane16_strm0_ready         ( DownstreamStackBusLane[17][16].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane16_strm0_cntl          ( DownstreamStackBusLane[17][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane16_strm0_data          ( DownstreamStackBusLane[17][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane16_strm0_data_valid    ( DownstreamStackBusLane[17][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane16_strm1_ready         ( DownstreamStackBusLane[17][16].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane16_strm1_cntl          ( DownstreamStackBusLane[17][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane16_strm1_data          ( DownstreamStackBusLane[17][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane16_strm1_data_valid    ( DownstreamStackBusLane[17][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane17_strm0_ready         ( DownstreamStackBusLane[17][17].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane17_strm0_cntl          ( DownstreamStackBusLane[17][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane17_strm0_data          ( DownstreamStackBusLane[17][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane17_strm0_data_valid    ( DownstreamStackBusLane[17][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane17_strm1_ready         ( DownstreamStackBusLane[17][17].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane17_strm1_cntl          ( DownstreamStackBusLane[17][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane17_strm1_data          ( DownstreamStackBusLane[17][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane17_strm1_data_valid    ( DownstreamStackBusLane[17][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane18_strm0_ready         ( DownstreamStackBusLane[17][18].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane18_strm0_cntl          ( DownstreamStackBusLane[17][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane18_strm0_data          ( DownstreamStackBusLane[17][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane18_strm0_data_valid    ( DownstreamStackBusLane[17][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane18_strm1_ready         ( DownstreamStackBusLane[17][18].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane18_strm1_cntl          ( DownstreamStackBusLane[17][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane18_strm1_data          ( DownstreamStackBusLane[17][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane18_strm1_data_valid    ( DownstreamStackBusLane[17][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane19_strm0_ready         ( DownstreamStackBusLane[17][19].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane19_strm0_cntl          ( DownstreamStackBusLane[17][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane19_strm0_data          ( DownstreamStackBusLane[17][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane19_strm0_data_valid    ( DownstreamStackBusLane[17][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane19_strm1_ready         ( DownstreamStackBusLane[17][19].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane19_strm1_cntl          ( DownstreamStackBusLane[17][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane19_strm1_data          ( DownstreamStackBusLane[17][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane19_strm1_data_valid    ( DownstreamStackBusLane[17][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane20_strm0_ready         ( DownstreamStackBusLane[17][20].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane20_strm0_cntl          ( DownstreamStackBusLane[17][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane20_strm0_data          ( DownstreamStackBusLane[17][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane20_strm0_data_valid    ( DownstreamStackBusLane[17][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane20_strm1_ready         ( DownstreamStackBusLane[17][20].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane20_strm1_cntl          ( DownstreamStackBusLane[17][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane20_strm1_data          ( DownstreamStackBusLane[17][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane20_strm1_data_valid    ( DownstreamStackBusLane[17][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane21_strm0_ready         ( DownstreamStackBusLane[17][21].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane21_strm0_cntl          ( DownstreamStackBusLane[17][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane21_strm0_data          ( DownstreamStackBusLane[17][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane21_strm0_data_valid    ( DownstreamStackBusLane[17][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane21_strm1_ready         ( DownstreamStackBusLane[17][21].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane21_strm1_cntl          ( DownstreamStackBusLane[17][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane21_strm1_data          ( DownstreamStackBusLane[17][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane21_strm1_data_valid    ( DownstreamStackBusLane[17][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane22_strm0_ready         ( DownstreamStackBusLane[17][22].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane22_strm0_cntl          ( DownstreamStackBusLane[17][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane22_strm0_data          ( DownstreamStackBusLane[17][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane22_strm0_data_valid    ( DownstreamStackBusLane[17][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane22_strm1_ready         ( DownstreamStackBusLane[17][22].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane22_strm1_cntl          ( DownstreamStackBusLane[17][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane22_strm1_data          ( DownstreamStackBusLane[17][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane22_strm1_data_valid    ( DownstreamStackBusLane[17][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane23_strm0_ready         ( DownstreamStackBusLane[17][23].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane23_strm0_cntl          ( DownstreamStackBusLane[17][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane23_strm0_data          ( DownstreamStackBusLane[17][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane23_strm0_data_valid    ( DownstreamStackBusLane[17][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane23_strm1_ready         ( DownstreamStackBusLane[17][23].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane23_strm1_cntl          ( DownstreamStackBusLane[17][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane23_strm1_data          ( DownstreamStackBusLane[17][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane23_strm1_data_valid    ( DownstreamStackBusLane[17][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane24_strm0_ready         ( DownstreamStackBusLane[17][24].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane24_strm0_cntl          ( DownstreamStackBusLane[17][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane24_strm0_data          ( DownstreamStackBusLane[17][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane24_strm0_data_valid    ( DownstreamStackBusLane[17][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane24_strm1_ready         ( DownstreamStackBusLane[17][24].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane24_strm1_cntl          ( DownstreamStackBusLane[17][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane24_strm1_data          ( DownstreamStackBusLane[17][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane24_strm1_data_valid    ( DownstreamStackBusLane[17][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane25_strm0_ready         ( DownstreamStackBusLane[17][25].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane25_strm0_cntl          ( DownstreamStackBusLane[17][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane25_strm0_data          ( DownstreamStackBusLane[17][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane25_strm0_data_valid    ( DownstreamStackBusLane[17][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane25_strm1_ready         ( DownstreamStackBusLane[17][25].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane25_strm1_cntl          ( DownstreamStackBusLane[17][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane25_strm1_data          ( DownstreamStackBusLane[17][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane25_strm1_data_valid    ( DownstreamStackBusLane[17][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane26_strm0_ready         ( DownstreamStackBusLane[17][26].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane26_strm0_cntl          ( DownstreamStackBusLane[17][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane26_strm0_data          ( DownstreamStackBusLane[17][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane26_strm0_data_valid    ( DownstreamStackBusLane[17][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane26_strm1_ready         ( DownstreamStackBusLane[17][26].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane26_strm1_cntl          ( DownstreamStackBusLane[17][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane26_strm1_data          ( DownstreamStackBusLane[17][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane26_strm1_data_valid    ( DownstreamStackBusLane[17][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane27_strm0_ready         ( DownstreamStackBusLane[17][27].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane27_strm0_cntl          ( DownstreamStackBusLane[17][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane27_strm0_data          ( DownstreamStackBusLane[17][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane27_strm0_data_valid    ( DownstreamStackBusLane[17][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane27_strm1_ready         ( DownstreamStackBusLane[17][27].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane27_strm1_cntl          ( DownstreamStackBusLane[17][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane27_strm1_data          ( DownstreamStackBusLane[17][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane27_strm1_data_valid    ( DownstreamStackBusLane[17][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane28_strm0_ready         ( DownstreamStackBusLane[17][28].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane28_strm0_cntl          ( DownstreamStackBusLane[17][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane28_strm0_data          ( DownstreamStackBusLane[17][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane28_strm0_data_valid    ( DownstreamStackBusLane[17][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane28_strm1_ready         ( DownstreamStackBusLane[17][28].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane28_strm1_cntl          ( DownstreamStackBusLane[17][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane28_strm1_data          ( DownstreamStackBusLane[17][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane28_strm1_data_valid    ( DownstreamStackBusLane[17][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane29_strm0_ready         ( DownstreamStackBusLane[17][29].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane29_strm0_cntl          ( DownstreamStackBusLane[17][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane29_strm0_data          ( DownstreamStackBusLane[17][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane29_strm0_data_valid    ( DownstreamStackBusLane[17][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane29_strm1_ready         ( DownstreamStackBusLane[17][29].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane29_strm1_cntl          ( DownstreamStackBusLane[17][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane29_strm1_data          ( DownstreamStackBusLane[17][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane29_strm1_data_valid    ( DownstreamStackBusLane[17][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane30_strm0_ready         ( DownstreamStackBusLane[17][30].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane30_strm0_cntl          ( DownstreamStackBusLane[17][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane30_strm0_data          ( DownstreamStackBusLane[17][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane30_strm0_data_valid    ( DownstreamStackBusLane[17][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane30_strm1_ready         ( DownstreamStackBusLane[17][30].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane30_strm1_cntl          ( DownstreamStackBusLane[17][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane30_strm1_data          ( DownstreamStackBusLane[17][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane30_strm1_data_valid    ( DownstreamStackBusLane[17][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 17, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane31_strm0_ready         ( DownstreamStackBusLane[17][31].pe__std__lane_strm0_ready              ),      
        .std__pe17__lane31_strm0_cntl          ( DownstreamStackBusLane[17][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe17__lane31_strm0_data          ( DownstreamStackBusLane[17][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe17__lane31_strm0_data_valid    ( DownstreamStackBusLane[17][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__std__lane31_strm1_ready         ( DownstreamStackBusLane[17][31].pe__std__lane_strm1_ready              ),      
        .std__pe17__lane31_strm1_cntl          ( DownstreamStackBusLane[17][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe17__lane31_strm1_data          ( DownstreamStackBusLane[17][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe17__lane31_strm1_data_valid    ( DownstreamStackBusLane[17][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane0_strm0_ready         ( DownstreamStackBusLane[18][0].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane0_strm0_cntl          ( DownstreamStackBusLane[18][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane0_strm0_data          ( DownstreamStackBusLane[18][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane0_strm0_data_valid    ( DownstreamStackBusLane[18][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane0_strm1_ready         ( DownstreamStackBusLane[18][0].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane0_strm1_cntl          ( DownstreamStackBusLane[18][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane0_strm1_data          ( DownstreamStackBusLane[18][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane0_strm1_data_valid    ( DownstreamStackBusLane[18][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane1_strm0_ready         ( DownstreamStackBusLane[18][1].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane1_strm0_cntl          ( DownstreamStackBusLane[18][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane1_strm0_data          ( DownstreamStackBusLane[18][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane1_strm0_data_valid    ( DownstreamStackBusLane[18][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane1_strm1_ready         ( DownstreamStackBusLane[18][1].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane1_strm1_cntl          ( DownstreamStackBusLane[18][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane1_strm1_data          ( DownstreamStackBusLane[18][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane1_strm1_data_valid    ( DownstreamStackBusLane[18][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane2_strm0_ready         ( DownstreamStackBusLane[18][2].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane2_strm0_cntl          ( DownstreamStackBusLane[18][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane2_strm0_data          ( DownstreamStackBusLane[18][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane2_strm0_data_valid    ( DownstreamStackBusLane[18][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane2_strm1_ready         ( DownstreamStackBusLane[18][2].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane2_strm1_cntl          ( DownstreamStackBusLane[18][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane2_strm1_data          ( DownstreamStackBusLane[18][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane2_strm1_data_valid    ( DownstreamStackBusLane[18][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane3_strm0_ready         ( DownstreamStackBusLane[18][3].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane3_strm0_cntl          ( DownstreamStackBusLane[18][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane3_strm0_data          ( DownstreamStackBusLane[18][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane3_strm0_data_valid    ( DownstreamStackBusLane[18][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane3_strm1_ready         ( DownstreamStackBusLane[18][3].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane3_strm1_cntl          ( DownstreamStackBusLane[18][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane3_strm1_data          ( DownstreamStackBusLane[18][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane3_strm1_data_valid    ( DownstreamStackBusLane[18][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane4_strm0_ready         ( DownstreamStackBusLane[18][4].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane4_strm0_cntl          ( DownstreamStackBusLane[18][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane4_strm0_data          ( DownstreamStackBusLane[18][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane4_strm0_data_valid    ( DownstreamStackBusLane[18][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane4_strm1_ready         ( DownstreamStackBusLane[18][4].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane4_strm1_cntl          ( DownstreamStackBusLane[18][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane4_strm1_data          ( DownstreamStackBusLane[18][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane4_strm1_data_valid    ( DownstreamStackBusLane[18][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane5_strm0_ready         ( DownstreamStackBusLane[18][5].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane5_strm0_cntl          ( DownstreamStackBusLane[18][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane5_strm0_data          ( DownstreamStackBusLane[18][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane5_strm0_data_valid    ( DownstreamStackBusLane[18][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane5_strm1_ready         ( DownstreamStackBusLane[18][5].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane5_strm1_cntl          ( DownstreamStackBusLane[18][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane5_strm1_data          ( DownstreamStackBusLane[18][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane5_strm1_data_valid    ( DownstreamStackBusLane[18][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane6_strm0_ready         ( DownstreamStackBusLane[18][6].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane6_strm0_cntl          ( DownstreamStackBusLane[18][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane6_strm0_data          ( DownstreamStackBusLane[18][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane6_strm0_data_valid    ( DownstreamStackBusLane[18][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane6_strm1_ready         ( DownstreamStackBusLane[18][6].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane6_strm1_cntl          ( DownstreamStackBusLane[18][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane6_strm1_data          ( DownstreamStackBusLane[18][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane6_strm1_data_valid    ( DownstreamStackBusLane[18][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane7_strm0_ready         ( DownstreamStackBusLane[18][7].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane7_strm0_cntl          ( DownstreamStackBusLane[18][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane7_strm0_data          ( DownstreamStackBusLane[18][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane7_strm0_data_valid    ( DownstreamStackBusLane[18][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane7_strm1_ready         ( DownstreamStackBusLane[18][7].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane7_strm1_cntl          ( DownstreamStackBusLane[18][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane7_strm1_data          ( DownstreamStackBusLane[18][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane7_strm1_data_valid    ( DownstreamStackBusLane[18][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane8_strm0_ready         ( DownstreamStackBusLane[18][8].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane8_strm0_cntl          ( DownstreamStackBusLane[18][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane8_strm0_data          ( DownstreamStackBusLane[18][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane8_strm0_data_valid    ( DownstreamStackBusLane[18][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane8_strm1_ready         ( DownstreamStackBusLane[18][8].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane8_strm1_cntl          ( DownstreamStackBusLane[18][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane8_strm1_data          ( DownstreamStackBusLane[18][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane8_strm1_data_valid    ( DownstreamStackBusLane[18][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane9_strm0_ready         ( DownstreamStackBusLane[18][9].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane9_strm0_cntl          ( DownstreamStackBusLane[18][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane9_strm0_data          ( DownstreamStackBusLane[18][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane9_strm0_data_valid    ( DownstreamStackBusLane[18][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane9_strm1_ready         ( DownstreamStackBusLane[18][9].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane9_strm1_cntl          ( DownstreamStackBusLane[18][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane9_strm1_data          ( DownstreamStackBusLane[18][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane9_strm1_data_valid    ( DownstreamStackBusLane[18][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane10_strm0_ready         ( DownstreamStackBusLane[18][10].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane10_strm0_cntl          ( DownstreamStackBusLane[18][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane10_strm0_data          ( DownstreamStackBusLane[18][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane10_strm0_data_valid    ( DownstreamStackBusLane[18][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane10_strm1_ready         ( DownstreamStackBusLane[18][10].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane10_strm1_cntl          ( DownstreamStackBusLane[18][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane10_strm1_data          ( DownstreamStackBusLane[18][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane10_strm1_data_valid    ( DownstreamStackBusLane[18][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane11_strm0_ready         ( DownstreamStackBusLane[18][11].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane11_strm0_cntl          ( DownstreamStackBusLane[18][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane11_strm0_data          ( DownstreamStackBusLane[18][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane11_strm0_data_valid    ( DownstreamStackBusLane[18][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane11_strm1_ready         ( DownstreamStackBusLane[18][11].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane11_strm1_cntl          ( DownstreamStackBusLane[18][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane11_strm1_data          ( DownstreamStackBusLane[18][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane11_strm1_data_valid    ( DownstreamStackBusLane[18][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane12_strm0_ready         ( DownstreamStackBusLane[18][12].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane12_strm0_cntl          ( DownstreamStackBusLane[18][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane12_strm0_data          ( DownstreamStackBusLane[18][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane12_strm0_data_valid    ( DownstreamStackBusLane[18][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane12_strm1_ready         ( DownstreamStackBusLane[18][12].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane12_strm1_cntl          ( DownstreamStackBusLane[18][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane12_strm1_data          ( DownstreamStackBusLane[18][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane12_strm1_data_valid    ( DownstreamStackBusLane[18][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane13_strm0_ready         ( DownstreamStackBusLane[18][13].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane13_strm0_cntl          ( DownstreamStackBusLane[18][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane13_strm0_data          ( DownstreamStackBusLane[18][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane13_strm0_data_valid    ( DownstreamStackBusLane[18][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane13_strm1_ready         ( DownstreamStackBusLane[18][13].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane13_strm1_cntl          ( DownstreamStackBusLane[18][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane13_strm1_data          ( DownstreamStackBusLane[18][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane13_strm1_data_valid    ( DownstreamStackBusLane[18][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane14_strm0_ready         ( DownstreamStackBusLane[18][14].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane14_strm0_cntl          ( DownstreamStackBusLane[18][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane14_strm0_data          ( DownstreamStackBusLane[18][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane14_strm0_data_valid    ( DownstreamStackBusLane[18][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane14_strm1_ready         ( DownstreamStackBusLane[18][14].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane14_strm1_cntl          ( DownstreamStackBusLane[18][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane14_strm1_data          ( DownstreamStackBusLane[18][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane14_strm1_data_valid    ( DownstreamStackBusLane[18][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane15_strm0_ready         ( DownstreamStackBusLane[18][15].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane15_strm0_cntl          ( DownstreamStackBusLane[18][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane15_strm0_data          ( DownstreamStackBusLane[18][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane15_strm0_data_valid    ( DownstreamStackBusLane[18][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane15_strm1_ready         ( DownstreamStackBusLane[18][15].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane15_strm1_cntl          ( DownstreamStackBusLane[18][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane15_strm1_data          ( DownstreamStackBusLane[18][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane15_strm1_data_valid    ( DownstreamStackBusLane[18][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane16_strm0_ready         ( DownstreamStackBusLane[18][16].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane16_strm0_cntl          ( DownstreamStackBusLane[18][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane16_strm0_data          ( DownstreamStackBusLane[18][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane16_strm0_data_valid    ( DownstreamStackBusLane[18][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane16_strm1_ready         ( DownstreamStackBusLane[18][16].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane16_strm1_cntl          ( DownstreamStackBusLane[18][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane16_strm1_data          ( DownstreamStackBusLane[18][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane16_strm1_data_valid    ( DownstreamStackBusLane[18][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane17_strm0_ready         ( DownstreamStackBusLane[18][17].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane17_strm0_cntl          ( DownstreamStackBusLane[18][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane17_strm0_data          ( DownstreamStackBusLane[18][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane17_strm0_data_valid    ( DownstreamStackBusLane[18][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane17_strm1_ready         ( DownstreamStackBusLane[18][17].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane17_strm1_cntl          ( DownstreamStackBusLane[18][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane17_strm1_data          ( DownstreamStackBusLane[18][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane17_strm1_data_valid    ( DownstreamStackBusLane[18][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane18_strm0_ready         ( DownstreamStackBusLane[18][18].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane18_strm0_cntl          ( DownstreamStackBusLane[18][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane18_strm0_data          ( DownstreamStackBusLane[18][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane18_strm0_data_valid    ( DownstreamStackBusLane[18][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane18_strm1_ready         ( DownstreamStackBusLane[18][18].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane18_strm1_cntl          ( DownstreamStackBusLane[18][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane18_strm1_data          ( DownstreamStackBusLane[18][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane18_strm1_data_valid    ( DownstreamStackBusLane[18][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane19_strm0_ready         ( DownstreamStackBusLane[18][19].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane19_strm0_cntl          ( DownstreamStackBusLane[18][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane19_strm0_data          ( DownstreamStackBusLane[18][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane19_strm0_data_valid    ( DownstreamStackBusLane[18][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane19_strm1_ready         ( DownstreamStackBusLane[18][19].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane19_strm1_cntl          ( DownstreamStackBusLane[18][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane19_strm1_data          ( DownstreamStackBusLane[18][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane19_strm1_data_valid    ( DownstreamStackBusLane[18][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane20_strm0_ready         ( DownstreamStackBusLane[18][20].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane20_strm0_cntl          ( DownstreamStackBusLane[18][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane20_strm0_data          ( DownstreamStackBusLane[18][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane20_strm0_data_valid    ( DownstreamStackBusLane[18][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane20_strm1_ready         ( DownstreamStackBusLane[18][20].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane20_strm1_cntl          ( DownstreamStackBusLane[18][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane20_strm1_data          ( DownstreamStackBusLane[18][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane20_strm1_data_valid    ( DownstreamStackBusLane[18][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane21_strm0_ready         ( DownstreamStackBusLane[18][21].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane21_strm0_cntl          ( DownstreamStackBusLane[18][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane21_strm0_data          ( DownstreamStackBusLane[18][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane21_strm0_data_valid    ( DownstreamStackBusLane[18][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane21_strm1_ready         ( DownstreamStackBusLane[18][21].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane21_strm1_cntl          ( DownstreamStackBusLane[18][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane21_strm1_data          ( DownstreamStackBusLane[18][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane21_strm1_data_valid    ( DownstreamStackBusLane[18][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane22_strm0_ready         ( DownstreamStackBusLane[18][22].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane22_strm0_cntl          ( DownstreamStackBusLane[18][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane22_strm0_data          ( DownstreamStackBusLane[18][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane22_strm0_data_valid    ( DownstreamStackBusLane[18][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane22_strm1_ready         ( DownstreamStackBusLane[18][22].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane22_strm1_cntl          ( DownstreamStackBusLane[18][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane22_strm1_data          ( DownstreamStackBusLane[18][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane22_strm1_data_valid    ( DownstreamStackBusLane[18][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane23_strm0_ready         ( DownstreamStackBusLane[18][23].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane23_strm0_cntl          ( DownstreamStackBusLane[18][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane23_strm0_data          ( DownstreamStackBusLane[18][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane23_strm0_data_valid    ( DownstreamStackBusLane[18][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane23_strm1_ready         ( DownstreamStackBusLane[18][23].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane23_strm1_cntl          ( DownstreamStackBusLane[18][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane23_strm1_data          ( DownstreamStackBusLane[18][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane23_strm1_data_valid    ( DownstreamStackBusLane[18][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane24_strm0_ready         ( DownstreamStackBusLane[18][24].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane24_strm0_cntl          ( DownstreamStackBusLane[18][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane24_strm0_data          ( DownstreamStackBusLane[18][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane24_strm0_data_valid    ( DownstreamStackBusLane[18][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane24_strm1_ready         ( DownstreamStackBusLane[18][24].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane24_strm1_cntl          ( DownstreamStackBusLane[18][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane24_strm1_data          ( DownstreamStackBusLane[18][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane24_strm1_data_valid    ( DownstreamStackBusLane[18][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane25_strm0_ready         ( DownstreamStackBusLane[18][25].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane25_strm0_cntl          ( DownstreamStackBusLane[18][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane25_strm0_data          ( DownstreamStackBusLane[18][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane25_strm0_data_valid    ( DownstreamStackBusLane[18][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane25_strm1_ready         ( DownstreamStackBusLane[18][25].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane25_strm1_cntl          ( DownstreamStackBusLane[18][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane25_strm1_data          ( DownstreamStackBusLane[18][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane25_strm1_data_valid    ( DownstreamStackBusLane[18][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane26_strm0_ready         ( DownstreamStackBusLane[18][26].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane26_strm0_cntl          ( DownstreamStackBusLane[18][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane26_strm0_data          ( DownstreamStackBusLane[18][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane26_strm0_data_valid    ( DownstreamStackBusLane[18][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane26_strm1_ready         ( DownstreamStackBusLane[18][26].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane26_strm1_cntl          ( DownstreamStackBusLane[18][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane26_strm1_data          ( DownstreamStackBusLane[18][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane26_strm1_data_valid    ( DownstreamStackBusLane[18][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane27_strm0_ready         ( DownstreamStackBusLane[18][27].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane27_strm0_cntl          ( DownstreamStackBusLane[18][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane27_strm0_data          ( DownstreamStackBusLane[18][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane27_strm0_data_valid    ( DownstreamStackBusLane[18][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane27_strm1_ready         ( DownstreamStackBusLane[18][27].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane27_strm1_cntl          ( DownstreamStackBusLane[18][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane27_strm1_data          ( DownstreamStackBusLane[18][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane27_strm1_data_valid    ( DownstreamStackBusLane[18][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane28_strm0_ready         ( DownstreamStackBusLane[18][28].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane28_strm0_cntl          ( DownstreamStackBusLane[18][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane28_strm0_data          ( DownstreamStackBusLane[18][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane28_strm0_data_valid    ( DownstreamStackBusLane[18][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane28_strm1_ready         ( DownstreamStackBusLane[18][28].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane28_strm1_cntl          ( DownstreamStackBusLane[18][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane28_strm1_data          ( DownstreamStackBusLane[18][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane28_strm1_data_valid    ( DownstreamStackBusLane[18][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane29_strm0_ready         ( DownstreamStackBusLane[18][29].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane29_strm0_cntl          ( DownstreamStackBusLane[18][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane29_strm0_data          ( DownstreamStackBusLane[18][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane29_strm0_data_valid    ( DownstreamStackBusLane[18][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane29_strm1_ready         ( DownstreamStackBusLane[18][29].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane29_strm1_cntl          ( DownstreamStackBusLane[18][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane29_strm1_data          ( DownstreamStackBusLane[18][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane29_strm1_data_valid    ( DownstreamStackBusLane[18][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane30_strm0_ready         ( DownstreamStackBusLane[18][30].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane30_strm0_cntl          ( DownstreamStackBusLane[18][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane30_strm0_data          ( DownstreamStackBusLane[18][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane30_strm0_data_valid    ( DownstreamStackBusLane[18][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane30_strm1_ready         ( DownstreamStackBusLane[18][30].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane30_strm1_cntl          ( DownstreamStackBusLane[18][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane30_strm1_data          ( DownstreamStackBusLane[18][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane30_strm1_data_valid    ( DownstreamStackBusLane[18][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 18, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane31_strm0_ready         ( DownstreamStackBusLane[18][31].pe__std__lane_strm0_ready              ),      
        .std__pe18__lane31_strm0_cntl          ( DownstreamStackBusLane[18][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe18__lane31_strm0_data          ( DownstreamStackBusLane[18][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe18__lane31_strm0_data_valid    ( DownstreamStackBusLane[18][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__std__lane31_strm1_ready         ( DownstreamStackBusLane[18][31].pe__std__lane_strm1_ready              ),      
        .std__pe18__lane31_strm1_cntl          ( DownstreamStackBusLane[18][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe18__lane31_strm1_data          ( DownstreamStackBusLane[18][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe18__lane31_strm1_data_valid    ( DownstreamStackBusLane[18][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane0_strm0_ready         ( DownstreamStackBusLane[19][0].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane0_strm0_cntl          ( DownstreamStackBusLane[19][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane0_strm0_data          ( DownstreamStackBusLane[19][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane0_strm0_data_valid    ( DownstreamStackBusLane[19][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane0_strm1_ready         ( DownstreamStackBusLane[19][0].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane0_strm1_cntl          ( DownstreamStackBusLane[19][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane0_strm1_data          ( DownstreamStackBusLane[19][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane0_strm1_data_valid    ( DownstreamStackBusLane[19][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane1_strm0_ready         ( DownstreamStackBusLane[19][1].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane1_strm0_cntl          ( DownstreamStackBusLane[19][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane1_strm0_data          ( DownstreamStackBusLane[19][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane1_strm0_data_valid    ( DownstreamStackBusLane[19][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane1_strm1_ready         ( DownstreamStackBusLane[19][1].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane1_strm1_cntl          ( DownstreamStackBusLane[19][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane1_strm1_data          ( DownstreamStackBusLane[19][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane1_strm1_data_valid    ( DownstreamStackBusLane[19][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane2_strm0_ready         ( DownstreamStackBusLane[19][2].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane2_strm0_cntl          ( DownstreamStackBusLane[19][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane2_strm0_data          ( DownstreamStackBusLane[19][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane2_strm0_data_valid    ( DownstreamStackBusLane[19][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane2_strm1_ready         ( DownstreamStackBusLane[19][2].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane2_strm1_cntl          ( DownstreamStackBusLane[19][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane2_strm1_data          ( DownstreamStackBusLane[19][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane2_strm1_data_valid    ( DownstreamStackBusLane[19][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane3_strm0_ready         ( DownstreamStackBusLane[19][3].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane3_strm0_cntl          ( DownstreamStackBusLane[19][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane3_strm0_data          ( DownstreamStackBusLane[19][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane3_strm0_data_valid    ( DownstreamStackBusLane[19][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane3_strm1_ready         ( DownstreamStackBusLane[19][3].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane3_strm1_cntl          ( DownstreamStackBusLane[19][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane3_strm1_data          ( DownstreamStackBusLane[19][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane3_strm1_data_valid    ( DownstreamStackBusLane[19][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane4_strm0_ready         ( DownstreamStackBusLane[19][4].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane4_strm0_cntl          ( DownstreamStackBusLane[19][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane4_strm0_data          ( DownstreamStackBusLane[19][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane4_strm0_data_valid    ( DownstreamStackBusLane[19][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane4_strm1_ready         ( DownstreamStackBusLane[19][4].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane4_strm1_cntl          ( DownstreamStackBusLane[19][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane4_strm1_data          ( DownstreamStackBusLane[19][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane4_strm1_data_valid    ( DownstreamStackBusLane[19][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane5_strm0_ready         ( DownstreamStackBusLane[19][5].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane5_strm0_cntl          ( DownstreamStackBusLane[19][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane5_strm0_data          ( DownstreamStackBusLane[19][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane5_strm0_data_valid    ( DownstreamStackBusLane[19][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane5_strm1_ready         ( DownstreamStackBusLane[19][5].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane5_strm1_cntl          ( DownstreamStackBusLane[19][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane5_strm1_data          ( DownstreamStackBusLane[19][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane5_strm1_data_valid    ( DownstreamStackBusLane[19][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane6_strm0_ready         ( DownstreamStackBusLane[19][6].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane6_strm0_cntl          ( DownstreamStackBusLane[19][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane6_strm0_data          ( DownstreamStackBusLane[19][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane6_strm0_data_valid    ( DownstreamStackBusLane[19][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane6_strm1_ready         ( DownstreamStackBusLane[19][6].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane6_strm1_cntl          ( DownstreamStackBusLane[19][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane6_strm1_data          ( DownstreamStackBusLane[19][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane6_strm1_data_valid    ( DownstreamStackBusLane[19][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane7_strm0_ready         ( DownstreamStackBusLane[19][7].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane7_strm0_cntl          ( DownstreamStackBusLane[19][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane7_strm0_data          ( DownstreamStackBusLane[19][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane7_strm0_data_valid    ( DownstreamStackBusLane[19][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane7_strm1_ready         ( DownstreamStackBusLane[19][7].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane7_strm1_cntl          ( DownstreamStackBusLane[19][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane7_strm1_data          ( DownstreamStackBusLane[19][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane7_strm1_data_valid    ( DownstreamStackBusLane[19][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane8_strm0_ready         ( DownstreamStackBusLane[19][8].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane8_strm0_cntl          ( DownstreamStackBusLane[19][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane8_strm0_data          ( DownstreamStackBusLane[19][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane8_strm0_data_valid    ( DownstreamStackBusLane[19][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane8_strm1_ready         ( DownstreamStackBusLane[19][8].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane8_strm1_cntl          ( DownstreamStackBusLane[19][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane8_strm1_data          ( DownstreamStackBusLane[19][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane8_strm1_data_valid    ( DownstreamStackBusLane[19][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane9_strm0_ready         ( DownstreamStackBusLane[19][9].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane9_strm0_cntl          ( DownstreamStackBusLane[19][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane9_strm0_data          ( DownstreamStackBusLane[19][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane9_strm0_data_valid    ( DownstreamStackBusLane[19][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane9_strm1_ready         ( DownstreamStackBusLane[19][9].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane9_strm1_cntl          ( DownstreamStackBusLane[19][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane9_strm1_data          ( DownstreamStackBusLane[19][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane9_strm1_data_valid    ( DownstreamStackBusLane[19][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane10_strm0_ready         ( DownstreamStackBusLane[19][10].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane10_strm0_cntl          ( DownstreamStackBusLane[19][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane10_strm0_data          ( DownstreamStackBusLane[19][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane10_strm0_data_valid    ( DownstreamStackBusLane[19][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane10_strm1_ready         ( DownstreamStackBusLane[19][10].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane10_strm1_cntl          ( DownstreamStackBusLane[19][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane10_strm1_data          ( DownstreamStackBusLane[19][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane10_strm1_data_valid    ( DownstreamStackBusLane[19][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane11_strm0_ready         ( DownstreamStackBusLane[19][11].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane11_strm0_cntl          ( DownstreamStackBusLane[19][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane11_strm0_data          ( DownstreamStackBusLane[19][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane11_strm0_data_valid    ( DownstreamStackBusLane[19][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane11_strm1_ready         ( DownstreamStackBusLane[19][11].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane11_strm1_cntl          ( DownstreamStackBusLane[19][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane11_strm1_data          ( DownstreamStackBusLane[19][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane11_strm1_data_valid    ( DownstreamStackBusLane[19][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane12_strm0_ready         ( DownstreamStackBusLane[19][12].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane12_strm0_cntl          ( DownstreamStackBusLane[19][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane12_strm0_data          ( DownstreamStackBusLane[19][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane12_strm0_data_valid    ( DownstreamStackBusLane[19][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane12_strm1_ready         ( DownstreamStackBusLane[19][12].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane12_strm1_cntl          ( DownstreamStackBusLane[19][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane12_strm1_data          ( DownstreamStackBusLane[19][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane12_strm1_data_valid    ( DownstreamStackBusLane[19][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane13_strm0_ready         ( DownstreamStackBusLane[19][13].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane13_strm0_cntl          ( DownstreamStackBusLane[19][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane13_strm0_data          ( DownstreamStackBusLane[19][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane13_strm0_data_valid    ( DownstreamStackBusLane[19][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane13_strm1_ready         ( DownstreamStackBusLane[19][13].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane13_strm1_cntl          ( DownstreamStackBusLane[19][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane13_strm1_data          ( DownstreamStackBusLane[19][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane13_strm1_data_valid    ( DownstreamStackBusLane[19][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane14_strm0_ready         ( DownstreamStackBusLane[19][14].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane14_strm0_cntl          ( DownstreamStackBusLane[19][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane14_strm0_data          ( DownstreamStackBusLane[19][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane14_strm0_data_valid    ( DownstreamStackBusLane[19][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane14_strm1_ready         ( DownstreamStackBusLane[19][14].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane14_strm1_cntl          ( DownstreamStackBusLane[19][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane14_strm1_data          ( DownstreamStackBusLane[19][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane14_strm1_data_valid    ( DownstreamStackBusLane[19][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane15_strm0_ready         ( DownstreamStackBusLane[19][15].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane15_strm0_cntl          ( DownstreamStackBusLane[19][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane15_strm0_data          ( DownstreamStackBusLane[19][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane15_strm0_data_valid    ( DownstreamStackBusLane[19][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane15_strm1_ready         ( DownstreamStackBusLane[19][15].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane15_strm1_cntl          ( DownstreamStackBusLane[19][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane15_strm1_data          ( DownstreamStackBusLane[19][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane15_strm1_data_valid    ( DownstreamStackBusLane[19][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane16_strm0_ready         ( DownstreamStackBusLane[19][16].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane16_strm0_cntl          ( DownstreamStackBusLane[19][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane16_strm0_data          ( DownstreamStackBusLane[19][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane16_strm0_data_valid    ( DownstreamStackBusLane[19][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane16_strm1_ready         ( DownstreamStackBusLane[19][16].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane16_strm1_cntl          ( DownstreamStackBusLane[19][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane16_strm1_data          ( DownstreamStackBusLane[19][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane16_strm1_data_valid    ( DownstreamStackBusLane[19][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane17_strm0_ready         ( DownstreamStackBusLane[19][17].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane17_strm0_cntl          ( DownstreamStackBusLane[19][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane17_strm0_data          ( DownstreamStackBusLane[19][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane17_strm0_data_valid    ( DownstreamStackBusLane[19][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane17_strm1_ready         ( DownstreamStackBusLane[19][17].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane17_strm1_cntl          ( DownstreamStackBusLane[19][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane17_strm1_data          ( DownstreamStackBusLane[19][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane17_strm1_data_valid    ( DownstreamStackBusLane[19][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane18_strm0_ready         ( DownstreamStackBusLane[19][18].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane18_strm0_cntl          ( DownstreamStackBusLane[19][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane18_strm0_data          ( DownstreamStackBusLane[19][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane18_strm0_data_valid    ( DownstreamStackBusLane[19][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane18_strm1_ready         ( DownstreamStackBusLane[19][18].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane18_strm1_cntl          ( DownstreamStackBusLane[19][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane18_strm1_data          ( DownstreamStackBusLane[19][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane18_strm1_data_valid    ( DownstreamStackBusLane[19][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane19_strm0_ready         ( DownstreamStackBusLane[19][19].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane19_strm0_cntl          ( DownstreamStackBusLane[19][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane19_strm0_data          ( DownstreamStackBusLane[19][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane19_strm0_data_valid    ( DownstreamStackBusLane[19][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane19_strm1_ready         ( DownstreamStackBusLane[19][19].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane19_strm1_cntl          ( DownstreamStackBusLane[19][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane19_strm1_data          ( DownstreamStackBusLane[19][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane19_strm1_data_valid    ( DownstreamStackBusLane[19][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane20_strm0_ready         ( DownstreamStackBusLane[19][20].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane20_strm0_cntl          ( DownstreamStackBusLane[19][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane20_strm0_data          ( DownstreamStackBusLane[19][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane20_strm0_data_valid    ( DownstreamStackBusLane[19][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane20_strm1_ready         ( DownstreamStackBusLane[19][20].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane20_strm1_cntl          ( DownstreamStackBusLane[19][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane20_strm1_data          ( DownstreamStackBusLane[19][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane20_strm1_data_valid    ( DownstreamStackBusLane[19][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane21_strm0_ready         ( DownstreamStackBusLane[19][21].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane21_strm0_cntl          ( DownstreamStackBusLane[19][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane21_strm0_data          ( DownstreamStackBusLane[19][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane21_strm0_data_valid    ( DownstreamStackBusLane[19][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane21_strm1_ready         ( DownstreamStackBusLane[19][21].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane21_strm1_cntl          ( DownstreamStackBusLane[19][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane21_strm1_data          ( DownstreamStackBusLane[19][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane21_strm1_data_valid    ( DownstreamStackBusLane[19][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane22_strm0_ready         ( DownstreamStackBusLane[19][22].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane22_strm0_cntl          ( DownstreamStackBusLane[19][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane22_strm0_data          ( DownstreamStackBusLane[19][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane22_strm0_data_valid    ( DownstreamStackBusLane[19][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane22_strm1_ready         ( DownstreamStackBusLane[19][22].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane22_strm1_cntl          ( DownstreamStackBusLane[19][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane22_strm1_data          ( DownstreamStackBusLane[19][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane22_strm1_data_valid    ( DownstreamStackBusLane[19][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane23_strm0_ready         ( DownstreamStackBusLane[19][23].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane23_strm0_cntl          ( DownstreamStackBusLane[19][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane23_strm0_data          ( DownstreamStackBusLane[19][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane23_strm0_data_valid    ( DownstreamStackBusLane[19][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane23_strm1_ready         ( DownstreamStackBusLane[19][23].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane23_strm1_cntl          ( DownstreamStackBusLane[19][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane23_strm1_data          ( DownstreamStackBusLane[19][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane23_strm1_data_valid    ( DownstreamStackBusLane[19][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane24_strm0_ready         ( DownstreamStackBusLane[19][24].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane24_strm0_cntl          ( DownstreamStackBusLane[19][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane24_strm0_data          ( DownstreamStackBusLane[19][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane24_strm0_data_valid    ( DownstreamStackBusLane[19][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane24_strm1_ready         ( DownstreamStackBusLane[19][24].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane24_strm1_cntl          ( DownstreamStackBusLane[19][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane24_strm1_data          ( DownstreamStackBusLane[19][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane24_strm1_data_valid    ( DownstreamStackBusLane[19][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane25_strm0_ready         ( DownstreamStackBusLane[19][25].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane25_strm0_cntl          ( DownstreamStackBusLane[19][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane25_strm0_data          ( DownstreamStackBusLane[19][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane25_strm0_data_valid    ( DownstreamStackBusLane[19][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane25_strm1_ready         ( DownstreamStackBusLane[19][25].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane25_strm1_cntl          ( DownstreamStackBusLane[19][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane25_strm1_data          ( DownstreamStackBusLane[19][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane25_strm1_data_valid    ( DownstreamStackBusLane[19][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane26_strm0_ready         ( DownstreamStackBusLane[19][26].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane26_strm0_cntl          ( DownstreamStackBusLane[19][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane26_strm0_data          ( DownstreamStackBusLane[19][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane26_strm0_data_valid    ( DownstreamStackBusLane[19][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane26_strm1_ready         ( DownstreamStackBusLane[19][26].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane26_strm1_cntl          ( DownstreamStackBusLane[19][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane26_strm1_data          ( DownstreamStackBusLane[19][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane26_strm1_data_valid    ( DownstreamStackBusLane[19][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane27_strm0_ready         ( DownstreamStackBusLane[19][27].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane27_strm0_cntl          ( DownstreamStackBusLane[19][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane27_strm0_data          ( DownstreamStackBusLane[19][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane27_strm0_data_valid    ( DownstreamStackBusLane[19][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane27_strm1_ready         ( DownstreamStackBusLane[19][27].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane27_strm1_cntl          ( DownstreamStackBusLane[19][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane27_strm1_data          ( DownstreamStackBusLane[19][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane27_strm1_data_valid    ( DownstreamStackBusLane[19][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane28_strm0_ready         ( DownstreamStackBusLane[19][28].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane28_strm0_cntl          ( DownstreamStackBusLane[19][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane28_strm0_data          ( DownstreamStackBusLane[19][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane28_strm0_data_valid    ( DownstreamStackBusLane[19][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane28_strm1_ready         ( DownstreamStackBusLane[19][28].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane28_strm1_cntl          ( DownstreamStackBusLane[19][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane28_strm1_data          ( DownstreamStackBusLane[19][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane28_strm1_data_valid    ( DownstreamStackBusLane[19][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane29_strm0_ready         ( DownstreamStackBusLane[19][29].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane29_strm0_cntl          ( DownstreamStackBusLane[19][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane29_strm0_data          ( DownstreamStackBusLane[19][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane29_strm0_data_valid    ( DownstreamStackBusLane[19][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane29_strm1_ready         ( DownstreamStackBusLane[19][29].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane29_strm1_cntl          ( DownstreamStackBusLane[19][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane29_strm1_data          ( DownstreamStackBusLane[19][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane29_strm1_data_valid    ( DownstreamStackBusLane[19][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane30_strm0_ready         ( DownstreamStackBusLane[19][30].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane30_strm0_cntl          ( DownstreamStackBusLane[19][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane30_strm0_data          ( DownstreamStackBusLane[19][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane30_strm0_data_valid    ( DownstreamStackBusLane[19][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane30_strm1_ready         ( DownstreamStackBusLane[19][30].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane30_strm1_cntl          ( DownstreamStackBusLane[19][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane30_strm1_data          ( DownstreamStackBusLane[19][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane30_strm1_data_valid    ( DownstreamStackBusLane[19][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 19, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane31_strm0_ready         ( DownstreamStackBusLane[19][31].pe__std__lane_strm0_ready              ),      
        .std__pe19__lane31_strm0_cntl          ( DownstreamStackBusLane[19][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe19__lane31_strm0_data          ( DownstreamStackBusLane[19][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe19__lane31_strm0_data_valid    ( DownstreamStackBusLane[19][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__std__lane31_strm1_ready         ( DownstreamStackBusLane[19][31].pe__std__lane_strm1_ready              ),      
        .std__pe19__lane31_strm1_cntl          ( DownstreamStackBusLane[19][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe19__lane31_strm1_data          ( DownstreamStackBusLane[19][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe19__lane31_strm1_data_valid    ( DownstreamStackBusLane[19][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane0_strm0_ready         ( DownstreamStackBusLane[20][0].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane0_strm0_cntl          ( DownstreamStackBusLane[20][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane0_strm0_data          ( DownstreamStackBusLane[20][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane0_strm0_data_valid    ( DownstreamStackBusLane[20][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane0_strm1_ready         ( DownstreamStackBusLane[20][0].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane0_strm1_cntl          ( DownstreamStackBusLane[20][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane0_strm1_data          ( DownstreamStackBusLane[20][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane0_strm1_data_valid    ( DownstreamStackBusLane[20][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane1_strm0_ready         ( DownstreamStackBusLane[20][1].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane1_strm0_cntl          ( DownstreamStackBusLane[20][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane1_strm0_data          ( DownstreamStackBusLane[20][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane1_strm0_data_valid    ( DownstreamStackBusLane[20][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane1_strm1_ready         ( DownstreamStackBusLane[20][1].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane1_strm1_cntl          ( DownstreamStackBusLane[20][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane1_strm1_data          ( DownstreamStackBusLane[20][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane1_strm1_data_valid    ( DownstreamStackBusLane[20][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane2_strm0_ready         ( DownstreamStackBusLane[20][2].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane2_strm0_cntl          ( DownstreamStackBusLane[20][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane2_strm0_data          ( DownstreamStackBusLane[20][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane2_strm0_data_valid    ( DownstreamStackBusLane[20][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane2_strm1_ready         ( DownstreamStackBusLane[20][2].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane2_strm1_cntl          ( DownstreamStackBusLane[20][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane2_strm1_data          ( DownstreamStackBusLane[20][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane2_strm1_data_valid    ( DownstreamStackBusLane[20][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane3_strm0_ready         ( DownstreamStackBusLane[20][3].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane3_strm0_cntl          ( DownstreamStackBusLane[20][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane3_strm0_data          ( DownstreamStackBusLane[20][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane3_strm0_data_valid    ( DownstreamStackBusLane[20][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane3_strm1_ready         ( DownstreamStackBusLane[20][3].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane3_strm1_cntl          ( DownstreamStackBusLane[20][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane3_strm1_data          ( DownstreamStackBusLane[20][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane3_strm1_data_valid    ( DownstreamStackBusLane[20][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane4_strm0_ready         ( DownstreamStackBusLane[20][4].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane4_strm0_cntl          ( DownstreamStackBusLane[20][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane4_strm0_data          ( DownstreamStackBusLane[20][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane4_strm0_data_valid    ( DownstreamStackBusLane[20][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane4_strm1_ready         ( DownstreamStackBusLane[20][4].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane4_strm1_cntl          ( DownstreamStackBusLane[20][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane4_strm1_data          ( DownstreamStackBusLane[20][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane4_strm1_data_valid    ( DownstreamStackBusLane[20][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane5_strm0_ready         ( DownstreamStackBusLane[20][5].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane5_strm0_cntl          ( DownstreamStackBusLane[20][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane5_strm0_data          ( DownstreamStackBusLane[20][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane5_strm0_data_valid    ( DownstreamStackBusLane[20][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane5_strm1_ready         ( DownstreamStackBusLane[20][5].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane5_strm1_cntl          ( DownstreamStackBusLane[20][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane5_strm1_data          ( DownstreamStackBusLane[20][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane5_strm1_data_valid    ( DownstreamStackBusLane[20][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane6_strm0_ready         ( DownstreamStackBusLane[20][6].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane6_strm0_cntl          ( DownstreamStackBusLane[20][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane6_strm0_data          ( DownstreamStackBusLane[20][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane6_strm0_data_valid    ( DownstreamStackBusLane[20][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane6_strm1_ready         ( DownstreamStackBusLane[20][6].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane6_strm1_cntl          ( DownstreamStackBusLane[20][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane6_strm1_data          ( DownstreamStackBusLane[20][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane6_strm1_data_valid    ( DownstreamStackBusLane[20][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane7_strm0_ready         ( DownstreamStackBusLane[20][7].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane7_strm0_cntl          ( DownstreamStackBusLane[20][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane7_strm0_data          ( DownstreamStackBusLane[20][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane7_strm0_data_valid    ( DownstreamStackBusLane[20][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane7_strm1_ready         ( DownstreamStackBusLane[20][7].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane7_strm1_cntl          ( DownstreamStackBusLane[20][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane7_strm1_data          ( DownstreamStackBusLane[20][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane7_strm1_data_valid    ( DownstreamStackBusLane[20][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane8_strm0_ready         ( DownstreamStackBusLane[20][8].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane8_strm0_cntl          ( DownstreamStackBusLane[20][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane8_strm0_data          ( DownstreamStackBusLane[20][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane8_strm0_data_valid    ( DownstreamStackBusLane[20][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane8_strm1_ready         ( DownstreamStackBusLane[20][8].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane8_strm1_cntl          ( DownstreamStackBusLane[20][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane8_strm1_data          ( DownstreamStackBusLane[20][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane8_strm1_data_valid    ( DownstreamStackBusLane[20][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane9_strm0_ready         ( DownstreamStackBusLane[20][9].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane9_strm0_cntl          ( DownstreamStackBusLane[20][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane9_strm0_data          ( DownstreamStackBusLane[20][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane9_strm0_data_valid    ( DownstreamStackBusLane[20][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane9_strm1_ready         ( DownstreamStackBusLane[20][9].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane9_strm1_cntl          ( DownstreamStackBusLane[20][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane9_strm1_data          ( DownstreamStackBusLane[20][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane9_strm1_data_valid    ( DownstreamStackBusLane[20][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane10_strm0_ready         ( DownstreamStackBusLane[20][10].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane10_strm0_cntl          ( DownstreamStackBusLane[20][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane10_strm0_data          ( DownstreamStackBusLane[20][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane10_strm0_data_valid    ( DownstreamStackBusLane[20][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane10_strm1_ready         ( DownstreamStackBusLane[20][10].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane10_strm1_cntl          ( DownstreamStackBusLane[20][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane10_strm1_data          ( DownstreamStackBusLane[20][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane10_strm1_data_valid    ( DownstreamStackBusLane[20][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane11_strm0_ready         ( DownstreamStackBusLane[20][11].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane11_strm0_cntl          ( DownstreamStackBusLane[20][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane11_strm0_data          ( DownstreamStackBusLane[20][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane11_strm0_data_valid    ( DownstreamStackBusLane[20][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane11_strm1_ready         ( DownstreamStackBusLane[20][11].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane11_strm1_cntl          ( DownstreamStackBusLane[20][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane11_strm1_data          ( DownstreamStackBusLane[20][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane11_strm1_data_valid    ( DownstreamStackBusLane[20][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane12_strm0_ready         ( DownstreamStackBusLane[20][12].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane12_strm0_cntl          ( DownstreamStackBusLane[20][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane12_strm0_data          ( DownstreamStackBusLane[20][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane12_strm0_data_valid    ( DownstreamStackBusLane[20][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane12_strm1_ready         ( DownstreamStackBusLane[20][12].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane12_strm1_cntl          ( DownstreamStackBusLane[20][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane12_strm1_data          ( DownstreamStackBusLane[20][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane12_strm1_data_valid    ( DownstreamStackBusLane[20][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane13_strm0_ready         ( DownstreamStackBusLane[20][13].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane13_strm0_cntl          ( DownstreamStackBusLane[20][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane13_strm0_data          ( DownstreamStackBusLane[20][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane13_strm0_data_valid    ( DownstreamStackBusLane[20][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane13_strm1_ready         ( DownstreamStackBusLane[20][13].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane13_strm1_cntl          ( DownstreamStackBusLane[20][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane13_strm1_data          ( DownstreamStackBusLane[20][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane13_strm1_data_valid    ( DownstreamStackBusLane[20][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane14_strm0_ready         ( DownstreamStackBusLane[20][14].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane14_strm0_cntl          ( DownstreamStackBusLane[20][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane14_strm0_data          ( DownstreamStackBusLane[20][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane14_strm0_data_valid    ( DownstreamStackBusLane[20][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane14_strm1_ready         ( DownstreamStackBusLane[20][14].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane14_strm1_cntl          ( DownstreamStackBusLane[20][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane14_strm1_data          ( DownstreamStackBusLane[20][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane14_strm1_data_valid    ( DownstreamStackBusLane[20][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane15_strm0_ready         ( DownstreamStackBusLane[20][15].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane15_strm0_cntl          ( DownstreamStackBusLane[20][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane15_strm0_data          ( DownstreamStackBusLane[20][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane15_strm0_data_valid    ( DownstreamStackBusLane[20][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane15_strm1_ready         ( DownstreamStackBusLane[20][15].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane15_strm1_cntl          ( DownstreamStackBusLane[20][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane15_strm1_data          ( DownstreamStackBusLane[20][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane15_strm1_data_valid    ( DownstreamStackBusLane[20][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane16_strm0_ready         ( DownstreamStackBusLane[20][16].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane16_strm0_cntl          ( DownstreamStackBusLane[20][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane16_strm0_data          ( DownstreamStackBusLane[20][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane16_strm0_data_valid    ( DownstreamStackBusLane[20][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane16_strm1_ready         ( DownstreamStackBusLane[20][16].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane16_strm1_cntl          ( DownstreamStackBusLane[20][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane16_strm1_data          ( DownstreamStackBusLane[20][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane16_strm1_data_valid    ( DownstreamStackBusLane[20][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane17_strm0_ready         ( DownstreamStackBusLane[20][17].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane17_strm0_cntl          ( DownstreamStackBusLane[20][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane17_strm0_data          ( DownstreamStackBusLane[20][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane17_strm0_data_valid    ( DownstreamStackBusLane[20][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane17_strm1_ready         ( DownstreamStackBusLane[20][17].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane17_strm1_cntl          ( DownstreamStackBusLane[20][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane17_strm1_data          ( DownstreamStackBusLane[20][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane17_strm1_data_valid    ( DownstreamStackBusLane[20][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane18_strm0_ready         ( DownstreamStackBusLane[20][18].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane18_strm0_cntl          ( DownstreamStackBusLane[20][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane18_strm0_data          ( DownstreamStackBusLane[20][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane18_strm0_data_valid    ( DownstreamStackBusLane[20][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane18_strm1_ready         ( DownstreamStackBusLane[20][18].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane18_strm1_cntl          ( DownstreamStackBusLane[20][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane18_strm1_data          ( DownstreamStackBusLane[20][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane18_strm1_data_valid    ( DownstreamStackBusLane[20][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane19_strm0_ready         ( DownstreamStackBusLane[20][19].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane19_strm0_cntl          ( DownstreamStackBusLane[20][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane19_strm0_data          ( DownstreamStackBusLane[20][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane19_strm0_data_valid    ( DownstreamStackBusLane[20][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane19_strm1_ready         ( DownstreamStackBusLane[20][19].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane19_strm1_cntl          ( DownstreamStackBusLane[20][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane19_strm1_data          ( DownstreamStackBusLane[20][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane19_strm1_data_valid    ( DownstreamStackBusLane[20][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane20_strm0_ready         ( DownstreamStackBusLane[20][20].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane20_strm0_cntl          ( DownstreamStackBusLane[20][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane20_strm0_data          ( DownstreamStackBusLane[20][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane20_strm0_data_valid    ( DownstreamStackBusLane[20][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane20_strm1_ready         ( DownstreamStackBusLane[20][20].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane20_strm1_cntl          ( DownstreamStackBusLane[20][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane20_strm1_data          ( DownstreamStackBusLane[20][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane20_strm1_data_valid    ( DownstreamStackBusLane[20][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane21_strm0_ready         ( DownstreamStackBusLane[20][21].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane21_strm0_cntl          ( DownstreamStackBusLane[20][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane21_strm0_data          ( DownstreamStackBusLane[20][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane21_strm0_data_valid    ( DownstreamStackBusLane[20][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane21_strm1_ready         ( DownstreamStackBusLane[20][21].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane21_strm1_cntl          ( DownstreamStackBusLane[20][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane21_strm1_data          ( DownstreamStackBusLane[20][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane21_strm1_data_valid    ( DownstreamStackBusLane[20][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane22_strm0_ready         ( DownstreamStackBusLane[20][22].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane22_strm0_cntl          ( DownstreamStackBusLane[20][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane22_strm0_data          ( DownstreamStackBusLane[20][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane22_strm0_data_valid    ( DownstreamStackBusLane[20][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane22_strm1_ready         ( DownstreamStackBusLane[20][22].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane22_strm1_cntl          ( DownstreamStackBusLane[20][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane22_strm1_data          ( DownstreamStackBusLane[20][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane22_strm1_data_valid    ( DownstreamStackBusLane[20][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane23_strm0_ready         ( DownstreamStackBusLane[20][23].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane23_strm0_cntl          ( DownstreamStackBusLane[20][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane23_strm0_data          ( DownstreamStackBusLane[20][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane23_strm0_data_valid    ( DownstreamStackBusLane[20][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane23_strm1_ready         ( DownstreamStackBusLane[20][23].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane23_strm1_cntl          ( DownstreamStackBusLane[20][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane23_strm1_data          ( DownstreamStackBusLane[20][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane23_strm1_data_valid    ( DownstreamStackBusLane[20][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane24_strm0_ready         ( DownstreamStackBusLane[20][24].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane24_strm0_cntl          ( DownstreamStackBusLane[20][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane24_strm0_data          ( DownstreamStackBusLane[20][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane24_strm0_data_valid    ( DownstreamStackBusLane[20][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane24_strm1_ready         ( DownstreamStackBusLane[20][24].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane24_strm1_cntl          ( DownstreamStackBusLane[20][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane24_strm1_data          ( DownstreamStackBusLane[20][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane24_strm1_data_valid    ( DownstreamStackBusLane[20][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane25_strm0_ready         ( DownstreamStackBusLane[20][25].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane25_strm0_cntl          ( DownstreamStackBusLane[20][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane25_strm0_data          ( DownstreamStackBusLane[20][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane25_strm0_data_valid    ( DownstreamStackBusLane[20][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane25_strm1_ready         ( DownstreamStackBusLane[20][25].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane25_strm1_cntl          ( DownstreamStackBusLane[20][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane25_strm1_data          ( DownstreamStackBusLane[20][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane25_strm1_data_valid    ( DownstreamStackBusLane[20][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane26_strm0_ready         ( DownstreamStackBusLane[20][26].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane26_strm0_cntl          ( DownstreamStackBusLane[20][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane26_strm0_data          ( DownstreamStackBusLane[20][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane26_strm0_data_valid    ( DownstreamStackBusLane[20][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane26_strm1_ready         ( DownstreamStackBusLane[20][26].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane26_strm1_cntl          ( DownstreamStackBusLane[20][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane26_strm1_data          ( DownstreamStackBusLane[20][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane26_strm1_data_valid    ( DownstreamStackBusLane[20][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane27_strm0_ready         ( DownstreamStackBusLane[20][27].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane27_strm0_cntl          ( DownstreamStackBusLane[20][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane27_strm0_data          ( DownstreamStackBusLane[20][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane27_strm0_data_valid    ( DownstreamStackBusLane[20][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane27_strm1_ready         ( DownstreamStackBusLane[20][27].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane27_strm1_cntl          ( DownstreamStackBusLane[20][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane27_strm1_data          ( DownstreamStackBusLane[20][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane27_strm1_data_valid    ( DownstreamStackBusLane[20][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane28_strm0_ready         ( DownstreamStackBusLane[20][28].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane28_strm0_cntl          ( DownstreamStackBusLane[20][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane28_strm0_data          ( DownstreamStackBusLane[20][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane28_strm0_data_valid    ( DownstreamStackBusLane[20][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane28_strm1_ready         ( DownstreamStackBusLane[20][28].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane28_strm1_cntl          ( DownstreamStackBusLane[20][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane28_strm1_data          ( DownstreamStackBusLane[20][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane28_strm1_data_valid    ( DownstreamStackBusLane[20][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane29_strm0_ready         ( DownstreamStackBusLane[20][29].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane29_strm0_cntl          ( DownstreamStackBusLane[20][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane29_strm0_data          ( DownstreamStackBusLane[20][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane29_strm0_data_valid    ( DownstreamStackBusLane[20][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane29_strm1_ready         ( DownstreamStackBusLane[20][29].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane29_strm1_cntl          ( DownstreamStackBusLane[20][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane29_strm1_data          ( DownstreamStackBusLane[20][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane29_strm1_data_valid    ( DownstreamStackBusLane[20][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane30_strm0_ready         ( DownstreamStackBusLane[20][30].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane30_strm0_cntl          ( DownstreamStackBusLane[20][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane30_strm0_data          ( DownstreamStackBusLane[20][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane30_strm0_data_valid    ( DownstreamStackBusLane[20][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane30_strm1_ready         ( DownstreamStackBusLane[20][30].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane30_strm1_cntl          ( DownstreamStackBusLane[20][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane30_strm1_data          ( DownstreamStackBusLane[20][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane30_strm1_data_valid    ( DownstreamStackBusLane[20][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 20, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane31_strm0_ready         ( DownstreamStackBusLane[20][31].pe__std__lane_strm0_ready              ),      
        .std__pe20__lane31_strm0_cntl          ( DownstreamStackBusLane[20][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe20__lane31_strm0_data          ( DownstreamStackBusLane[20][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe20__lane31_strm0_data_valid    ( DownstreamStackBusLane[20][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__std__lane31_strm1_ready         ( DownstreamStackBusLane[20][31].pe__std__lane_strm1_ready              ),      
        .std__pe20__lane31_strm1_cntl          ( DownstreamStackBusLane[20][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe20__lane31_strm1_data          ( DownstreamStackBusLane[20][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe20__lane31_strm1_data_valid    ( DownstreamStackBusLane[20][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane0_strm0_ready         ( DownstreamStackBusLane[21][0].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane0_strm0_cntl          ( DownstreamStackBusLane[21][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane0_strm0_data          ( DownstreamStackBusLane[21][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane0_strm0_data_valid    ( DownstreamStackBusLane[21][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane0_strm1_ready         ( DownstreamStackBusLane[21][0].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane0_strm1_cntl          ( DownstreamStackBusLane[21][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane0_strm1_data          ( DownstreamStackBusLane[21][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane0_strm1_data_valid    ( DownstreamStackBusLane[21][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane1_strm0_ready         ( DownstreamStackBusLane[21][1].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane1_strm0_cntl          ( DownstreamStackBusLane[21][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane1_strm0_data          ( DownstreamStackBusLane[21][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane1_strm0_data_valid    ( DownstreamStackBusLane[21][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane1_strm1_ready         ( DownstreamStackBusLane[21][1].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane1_strm1_cntl          ( DownstreamStackBusLane[21][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane1_strm1_data          ( DownstreamStackBusLane[21][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane1_strm1_data_valid    ( DownstreamStackBusLane[21][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane2_strm0_ready         ( DownstreamStackBusLane[21][2].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane2_strm0_cntl          ( DownstreamStackBusLane[21][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane2_strm0_data          ( DownstreamStackBusLane[21][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane2_strm0_data_valid    ( DownstreamStackBusLane[21][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane2_strm1_ready         ( DownstreamStackBusLane[21][2].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane2_strm1_cntl          ( DownstreamStackBusLane[21][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane2_strm1_data          ( DownstreamStackBusLane[21][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane2_strm1_data_valid    ( DownstreamStackBusLane[21][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane3_strm0_ready         ( DownstreamStackBusLane[21][3].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane3_strm0_cntl          ( DownstreamStackBusLane[21][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane3_strm0_data          ( DownstreamStackBusLane[21][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane3_strm0_data_valid    ( DownstreamStackBusLane[21][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane3_strm1_ready         ( DownstreamStackBusLane[21][3].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane3_strm1_cntl          ( DownstreamStackBusLane[21][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane3_strm1_data          ( DownstreamStackBusLane[21][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane3_strm1_data_valid    ( DownstreamStackBusLane[21][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane4_strm0_ready         ( DownstreamStackBusLane[21][4].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane4_strm0_cntl          ( DownstreamStackBusLane[21][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane4_strm0_data          ( DownstreamStackBusLane[21][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane4_strm0_data_valid    ( DownstreamStackBusLane[21][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane4_strm1_ready         ( DownstreamStackBusLane[21][4].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane4_strm1_cntl          ( DownstreamStackBusLane[21][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane4_strm1_data          ( DownstreamStackBusLane[21][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane4_strm1_data_valid    ( DownstreamStackBusLane[21][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane5_strm0_ready         ( DownstreamStackBusLane[21][5].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane5_strm0_cntl          ( DownstreamStackBusLane[21][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane5_strm0_data          ( DownstreamStackBusLane[21][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane5_strm0_data_valid    ( DownstreamStackBusLane[21][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane5_strm1_ready         ( DownstreamStackBusLane[21][5].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane5_strm1_cntl          ( DownstreamStackBusLane[21][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane5_strm1_data          ( DownstreamStackBusLane[21][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane5_strm1_data_valid    ( DownstreamStackBusLane[21][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane6_strm0_ready         ( DownstreamStackBusLane[21][6].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane6_strm0_cntl          ( DownstreamStackBusLane[21][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane6_strm0_data          ( DownstreamStackBusLane[21][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane6_strm0_data_valid    ( DownstreamStackBusLane[21][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane6_strm1_ready         ( DownstreamStackBusLane[21][6].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane6_strm1_cntl          ( DownstreamStackBusLane[21][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane6_strm1_data          ( DownstreamStackBusLane[21][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane6_strm1_data_valid    ( DownstreamStackBusLane[21][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane7_strm0_ready         ( DownstreamStackBusLane[21][7].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane7_strm0_cntl          ( DownstreamStackBusLane[21][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane7_strm0_data          ( DownstreamStackBusLane[21][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane7_strm0_data_valid    ( DownstreamStackBusLane[21][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane7_strm1_ready         ( DownstreamStackBusLane[21][7].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane7_strm1_cntl          ( DownstreamStackBusLane[21][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane7_strm1_data          ( DownstreamStackBusLane[21][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane7_strm1_data_valid    ( DownstreamStackBusLane[21][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane8_strm0_ready         ( DownstreamStackBusLane[21][8].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane8_strm0_cntl          ( DownstreamStackBusLane[21][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane8_strm0_data          ( DownstreamStackBusLane[21][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane8_strm0_data_valid    ( DownstreamStackBusLane[21][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane8_strm1_ready         ( DownstreamStackBusLane[21][8].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane8_strm1_cntl          ( DownstreamStackBusLane[21][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane8_strm1_data          ( DownstreamStackBusLane[21][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane8_strm1_data_valid    ( DownstreamStackBusLane[21][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane9_strm0_ready         ( DownstreamStackBusLane[21][9].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane9_strm0_cntl          ( DownstreamStackBusLane[21][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane9_strm0_data          ( DownstreamStackBusLane[21][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane9_strm0_data_valid    ( DownstreamStackBusLane[21][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane9_strm1_ready         ( DownstreamStackBusLane[21][9].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane9_strm1_cntl          ( DownstreamStackBusLane[21][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane9_strm1_data          ( DownstreamStackBusLane[21][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane9_strm1_data_valid    ( DownstreamStackBusLane[21][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane10_strm0_ready         ( DownstreamStackBusLane[21][10].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane10_strm0_cntl          ( DownstreamStackBusLane[21][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane10_strm0_data          ( DownstreamStackBusLane[21][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane10_strm0_data_valid    ( DownstreamStackBusLane[21][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane10_strm1_ready         ( DownstreamStackBusLane[21][10].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane10_strm1_cntl          ( DownstreamStackBusLane[21][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane10_strm1_data          ( DownstreamStackBusLane[21][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane10_strm1_data_valid    ( DownstreamStackBusLane[21][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane11_strm0_ready         ( DownstreamStackBusLane[21][11].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane11_strm0_cntl          ( DownstreamStackBusLane[21][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane11_strm0_data          ( DownstreamStackBusLane[21][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane11_strm0_data_valid    ( DownstreamStackBusLane[21][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane11_strm1_ready         ( DownstreamStackBusLane[21][11].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane11_strm1_cntl          ( DownstreamStackBusLane[21][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane11_strm1_data          ( DownstreamStackBusLane[21][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane11_strm1_data_valid    ( DownstreamStackBusLane[21][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane12_strm0_ready         ( DownstreamStackBusLane[21][12].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane12_strm0_cntl          ( DownstreamStackBusLane[21][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane12_strm0_data          ( DownstreamStackBusLane[21][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane12_strm0_data_valid    ( DownstreamStackBusLane[21][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane12_strm1_ready         ( DownstreamStackBusLane[21][12].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane12_strm1_cntl          ( DownstreamStackBusLane[21][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane12_strm1_data          ( DownstreamStackBusLane[21][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane12_strm1_data_valid    ( DownstreamStackBusLane[21][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane13_strm0_ready         ( DownstreamStackBusLane[21][13].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane13_strm0_cntl          ( DownstreamStackBusLane[21][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane13_strm0_data          ( DownstreamStackBusLane[21][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane13_strm0_data_valid    ( DownstreamStackBusLane[21][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane13_strm1_ready         ( DownstreamStackBusLane[21][13].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane13_strm1_cntl          ( DownstreamStackBusLane[21][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane13_strm1_data          ( DownstreamStackBusLane[21][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane13_strm1_data_valid    ( DownstreamStackBusLane[21][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane14_strm0_ready         ( DownstreamStackBusLane[21][14].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane14_strm0_cntl          ( DownstreamStackBusLane[21][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane14_strm0_data          ( DownstreamStackBusLane[21][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane14_strm0_data_valid    ( DownstreamStackBusLane[21][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane14_strm1_ready         ( DownstreamStackBusLane[21][14].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane14_strm1_cntl          ( DownstreamStackBusLane[21][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane14_strm1_data          ( DownstreamStackBusLane[21][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane14_strm1_data_valid    ( DownstreamStackBusLane[21][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane15_strm0_ready         ( DownstreamStackBusLane[21][15].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane15_strm0_cntl          ( DownstreamStackBusLane[21][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane15_strm0_data          ( DownstreamStackBusLane[21][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane15_strm0_data_valid    ( DownstreamStackBusLane[21][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane15_strm1_ready         ( DownstreamStackBusLane[21][15].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane15_strm1_cntl          ( DownstreamStackBusLane[21][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane15_strm1_data          ( DownstreamStackBusLane[21][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane15_strm1_data_valid    ( DownstreamStackBusLane[21][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane16_strm0_ready         ( DownstreamStackBusLane[21][16].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane16_strm0_cntl          ( DownstreamStackBusLane[21][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane16_strm0_data          ( DownstreamStackBusLane[21][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane16_strm0_data_valid    ( DownstreamStackBusLane[21][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane16_strm1_ready         ( DownstreamStackBusLane[21][16].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane16_strm1_cntl          ( DownstreamStackBusLane[21][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane16_strm1_data          ( DownstreamStackBusLane[21][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane16_strm1_data_valid    ( DownstreamStackBusLane[21][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane17_strm0_ready         ( DownstreamStackBusLane[21][17].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane17_strm0_cntl          ( DownstreamStackBusLane[21][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane17_strm0_data          ( DownstreamStackBusLane[21][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane17_strm0_data_valid    ( DownstreamStackBusLane[21][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane17_strm1_ready         ( DownstreamStackBusLane[21][17].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane17_strm1_cntl          ( DownstreamStackBusLane[21][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane17_strm1_data          ( DownstreamStackBusLane[21][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane17_strm1_data_valid    ( DownstreamStackBusLane[21][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane18_strm0_ready         ( DownstreamStackBusLane[21][18].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane18_strm0_cntl          ( DownstreamStackBusLane[21][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane18_strm0_data          ( DownstreamStackBusLane[21][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane18_strm0_data_valid    ( DownstreamStackBusLane[21][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane18_strm1_ready         ( DownstreamStackBusLane[21][18].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane18_strm1_cntl          ( DownstreamStackBusLane[21][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane18_strm1_data          ( DownstreamStackBusLane[21][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane18_strm1_data_valid    ( DownstreamStackBusLane[21][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane19_strm0_ready         ( DownstreamStackBusLane[21][19].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane19_strm0_cntl          ( DownstreamStackBusLane[21][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane19_strm0_data          ( DownstreamStackBusLane[21][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane19_strm0_data_valid    ( DownstreamStackBusLane[21][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane19_strm1_ready         ( DownstreamStackBusLane[21][19].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane19_strm1_cntl          ( DownstreamStackBusLane[21][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane19_strm1_data          ( DownstreamStackBusLane[21][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane19_strm1_data_valid    ( DownstreamStackBusLane[21][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane20_strm0_ready         ( DownstreamStackBusLane[21][20].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane20_strm0_cntl          ( DownstreamStackBusLane[21][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane20_strm0_data          ( DownstreamStackBusLane[21][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane20_strm0_data_valid    ( DownstreamStackBusLane[21][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane20_strm1_ready         ( DownstreamStackBusLane[21][20].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane20_strm1_cntl          ( DownstreamStackBusLane[21][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane20_strm1_data          ( DownstreamStackBusLane[21][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane20_strm1_data_valid    ( DownstreamStackBusLane[21][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane21_strm0_ready         ( DownstreamStackBusLane[21][21].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane21_strm0_cntl          ( DownstreamStackBusLane[21][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane21_strm0_data          ( DownstreamStackBusLane[21][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane21_strm0_data_valid    ( DownstreamStackBusLane[21][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane21_strm1_ready         ( DownstreamStackBusLane[21][21].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane21_strm1_cntl          ( DownstreamStackBusLane[21][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane21_strm1_data          ( DownstreamStackBusLane[21][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane21_strm1_data_valid    ( DownstreamStackBusLane[21][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane22_strm0_ready         ( DownstreamStackBusLane[21][22].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane22_strm0_cntl          ( DownstreamStackBusLane[21][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane22_strm0_data          ( DownstreamStackBusLane[21][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane22_strm0_data_valid    ( DownstreamStackBusLane[21][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane22_strm1_ready         ( DownstreamStackBusLane[21][22].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane22_strm1_cntl          ( DownstreamStackBusLane[21][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane22_strm1_data          ( DownstreamStackBusLane[21][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane22_strm1_data_valid    ( DownstreamStackBusLane[21][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane23_strm0_ready         ( DownstreamStackBusLane[21][23].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane23_strm0_cntl          ( DownstreamStackBusLane[21][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane23_strm0_data          ( DownstreamStackBusLane[21][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane23_strm0_data_valid    ( DownstreamStackBusLane[21][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane23_strm1_ready         ( DownstreamStackBusLane[21][23].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane23_strm1_cntl          ( DownstreamStackBusLane[21][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane23_strm1_data          ( DownstreamStackBusLane[21][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane23_strm1_data_valid    ( DownstreamStackBusLane[21][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane24_strm0_ready         ( DownstreamStackBusLane[21][24].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane24_strm0_cntl          ( DownstreamStackBusLane[21][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane24_strm0_data          ( DownstreamStackBusLane[21][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane24_strm0_data_valid    ( DownstreamStackBusLane[21][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane24_strm1_ready         ( DownstreamStackBusLane[21][24].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane24_strm1_cntl          ( DownstreamStackBusLane[21][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane24_strm1_data          ( DownstreamStackBusLane[21][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane24_strm1_data_valid    ( DownstreamStackBusLane[21][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane25_strm0_ready         ( DownstreamStackBusLane[21][25].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane25_strm0_cntl          ( DownstreamStackBusLane[21][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane25_strm0_data          ( DownstreamStackBusLane[21][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane25_strm0_data_valid    ( DownstreamStackBusLane[21][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane25_strm1_ready         ( DownstreamStackBusLane[21][25].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane25_strm1_cntl          ( DownstreamStackBusLane[21][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane25_strm1_data          ( DownstreamStackBusLane[21][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane25_strm1_data_valid    ( DownstreamStackBusLane[21][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane26_strm0_ready         ( DownstreamStackBusLane[21][26].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane26_strm0_cntl          ( DownstreamStackBusLane[21][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane26_strm0_data          ( DownstreamStackBusLane[21][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane26_strm0_data_valid    ( DownstreamStackBusLane[21][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane26_strm1_ready         ( DownstreamStackBusLane[21][26].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane26_strm1_cntl          ( DownstreamStackBusLane[21][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane26_strm1_data          ( DownstreamStackBusLane[21][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane26_strm1_data_valid    ( DownstreamStackBusLane[21][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane27_strm0_ready         ( DownstreamStackBusLane[21][27].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane27_strm0_cntl          ( DownstreamStackBusLane[21][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane27_strm0_data          ( DownstreamStackBusLane[21][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane27_strm0_data_valid    ( DownstreamStackBusLane[21][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane27_strm1_ready         ( DownstreamStackBusLane[21][27].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane27_strm1_cntl          ( DownstreamStackBusLane[21][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane27_strm1_data          ( DownstreamStackBusLane[21][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane27_strm1_data_valid    ( DownstreamStackBusLane[21][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane28_strm0_ready         ( DownstreamStackBusLane[21][28].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane28_strm0_cntl          ( DownstreamStackBusLane[21][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane28_strm0_data          ( DownstreamStackBusLane[21][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane28_strm0_data_valid    ( DownstreamStackBusLane[21][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane28_strm1_ready         ( DownstreamStackBusLane[21][28].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane28_strm1_cntl          ( DownstreamStackBusLane[21][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane28_strm1_data          ( DownstreamStackBusLane[21][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane28_strm1_data_valid    ( DownstreamStackBusLane[21][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane29_strm0_ready         ( DownstreamStackBusLane[21][29].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane29_strm0_cntl          ( DownstreamStackBusLane[21][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane29_strm0_data          ( DownstreamStackBusLane[21][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane29_strm0_data_valid    ( DownstreamStackBusLane[21][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane29_strm1_ready         ( DownstreamStackBusLane[21][29].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane29_strm1_cntl          ( DownstreamStackBusLane[21][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane29_strm1_data          ( DownstreamStackBusLane[21][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane29_strm1_data_valid    ( DownstreamStackBusLane[21][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane30_strm0_ready         ( DownstreamStackBusLane[21][30].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane30_strm0_cntl          ( DownstreamStackBusLane[21][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane30_strm0_data          ( DownstreamStackBusLane[21][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane30_strm0_data_valid    ( DownstreamStackBusLane[21][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane30_strm1_ready         ( DownstreamStackBusLane[21][30].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane30_strm1_cntl          ( DownstreamStackBusLane[21][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane30_strm1_data          ( DownstreamStackBusLane[21][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane30_strm1_data_valid    ( DownstreamStackBusLane[21][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 21, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane31_strm0_ready         ( DownstreamStackBusLane[21][31].pe__std__lane_strm0_ready              ),      
        .std__pe21__lane31_strm0_cntl          ( DownstreamStackBusLane[21][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe21__lane31_strm0_data          ( DownstreamStackBusLane[21][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe21__lane31_strm0_data_valid    ( DownstreamStackBusLane[21][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__std__lane31_strm1_ready         ( DownstreamStackBusLane[21][31].pe__std__lane_strm1_ready              ),      
        .std__pe21__lane31_strm1_cntl          ( DownstreamStackBusLane[21][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe21__lane31_strm1_data          ( DownstreamStackBusLane[21][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe21__lane31_strm1_data_valid    ( DownstreamStackBusLane[21][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane0_strm0_ready         ( DownstreamStackBusLane[22][0].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane0_strm0_cntl          ( DownstreamStackBusLane[22][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane0_strm0_data          ( DownstreamStackBusLane[22][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane0_strm0_data_valid    ( DownstreamStackBusLane[22][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane0_strm1_ready         ( DownstreamStackBusLane[22][0].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane0_strm1_cntl          ( DownstreamStackBusLane[22][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane0_strm1_data          ( DownstreamStackBusLane[22][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane0_strm1_data_valid    ( DownstreamStackBusLane[22][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane1_strm0_ready         ( DownstreamStackBusLane[22][1].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane1_strm0_cntl          ( DownstreamStackBusLane[22][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane1_strm0_data          ( DownstreamStackBusLane[22][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane1_strm0_data_valid    ( DownstreamStackBusLane[22][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane1_strm1_ready         ( DownstreamStackBusLane[22][1].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane1_strm1_cntl          ( DownstreamStackBusLane[22][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane1_strm1_data          ( DownstreamStackBusLane[22][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane1_strm1_data_valid    ( DownstreamStackBusLane[22][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane2_strm0_ready         ( DownstreamStackBusLane[22][2].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane2_strm0_cntl          ( DownstreamStackBusLane[22][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane2_strm0_data          ( DownstreamStackBusLane[22][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane2_strm0_data_valid    ( DownstreamStackBusLane[22][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane2_strm1_ready         ( DownstreamStackBusLane[22][2].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane2_strm1_cntl          ( DownstreamStackBusLane[22][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane2_strm1_data          ( DownstreamStackBusLane[22][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane2_strm1_data_valid    ( DownstreamStackBusLane[22][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane3_strm0_ready         ( DownstreamStackBusLane[22][3].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane3_strm0_cntl          ( DownstreamStackBusLane[22][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane3_strm0_data          ( DownstreamStackBusLane[22][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane3_strm0_data_valid    ( DownstreamStackBusLane[22][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane3_strm1_ready         ( DownstreamStackBusLane[22][3].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane3_strm1_cntl          ( DownstreamStackBusLane[22][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane3_strm1_data          ( DownstreamStackBusLane[22][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane3_strm1_data_valid    ( DownstreamStackBusLane[22][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane4_strm0_ready         ( DownstreamStackBusLane[22][4].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane4_strm0_cntl          ( DownstreamStackBusLane[22][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane4_strm0_data          ( DownstreamStackBusLane[22][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane4_strm0_data_valid    ( DownstreamStackBusLane[22][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane4_strm1_ready         ( DownstreamStackBusLane[22][4].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane4_strm1_cntl          ( DownstreamStackBusLane[22][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane4_strm1_data          ( DownstreamStackBusLane[22][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane4_strm1_data_valid    ( DownstreamStackBusLane[22][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane5_strm0_ready         ( DownstreamStackBusLane[22][5].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane5_strm0_cntl          ( DownstreamStackBusLane[22][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane5_strm0_data          ( DownstreamStackBusLane[22][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane5_strm0_data_valid    ( DownstreamStackBusLane[22][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane5_strm1_ready         ( DownstreamStackBusLane[22][5].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane5_strm1_cntl          ( DownstreamStackBusLane[22][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane5_strm1_data          ( DownstreamStackBusLane[22][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane5_strm1_data_valid    ( DownstreamStackBusLane[22][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane6_strm0_ready         ( DownstreamStackBusLane[22][6].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane6_strm0_cntl          ( DownstreamStackBusLane[22][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane6_strm0_data          ( DownstreamStackBusLane[22][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane6_strm0_data_valid    ( DownstreamStackBusLane[22][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane6_strm1_ready         ( DownstreamStackBusLane[22][6].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane6_strm1_cntl          ( DownstreamStackBusLane[22][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane6_strm1_data          ( DownstreamStackBusLane[22][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane6_strm1_data_valid    ( DownstreamStackBusLane[22][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane7_strm0_ready         ( DownstreamStackBusLane[22][7].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane7_strm0_cntl          ( DownstreamStackBusLane[22][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane7_strm0_data          ( DownstreamStackBusLane[22][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane7_strm0_data_valid    ( DownstreamStackBusLane[22][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane7_strm1_ready         ( DownstreamStackBusLane[22][7].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane7_strm1_cntl          ( DownstreamStackBusLane[22][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane7_strm1_data          ( DownstreamStackBusLane[22][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane7_strm1_data_valid    ( DownstreamStackBusLane[22][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane8_strm0_ready         ( DownstreamStackBusLane[22][8].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane8_strm0_cntl          ( DownstreamStackBusLane[22][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane8_strm0_data          ( DownstreamStackBusLane[22][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane8_strm0_data_valid    ( DownstreamStackBusLane[22][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane8_strm1_ready         ( DownstreamStackBusLane[22][8].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane8_strm1_cntl          ( DownstreamStackBusLane[22][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane8_strm1_data          ( DownstreamStackBusLane[22][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane8_strm1_data_valid    ( DownstreamStackBusLane[22][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane9_strm0_ready         ( DownstreamStackBusLane[22][9].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane9_strm0_cntl          ( DownstreamStackBusLane[22][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane9_strm0_data          ( DownstreamStackBusLane[22][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane9_strm0_data_valid    ( DownstreamStackBusLane[22][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane9_strm1_ready         ( DownstreamStackBusLane[22][9].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane9_strm1_cntl          ( DownstreamStackBusLane[22][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane9_strm1_data          ( DownstreamStackBusLane[22][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane9_strm1_data_valid    ( DownstreamStackBusLane[22][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane10_strm0_ready         ( DownstreamStackBusLane[22][10].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane10_strm0_cntl          ( DownstreamStackBusLane[22][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane10_strm0_data          ( DownstreamStackBusLane[22][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane10_strm0_data_valid    ( DownstreamStackBusLane[22][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane10_strm1_ready         ( DownstreamStackBusLane[22][10].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane10_strm1_cntl          ( DownstreamStackBusLane[22][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane10_strm1_data          ( DownstreamStackBusLane[22][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane10_strm1_data_valid    ( DownstreamStackBusLane[22][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane11_strm0_ready         ( DownstreamStackBusLane[22][11].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane11_strm0_cntl          ( DownstreamStackBusLane[22][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane11_strm0_data          ( DownstreamStackBusLane[22][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane11_strm0_data_valid    ( DownstreamStackBusLane[22][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane11_strm1_ready         ( DownstreamStackBusLane[22][11].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane11_strm1_cntl          ( DownstreamStackBusLane[22][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane11_strm1_data          ( DownstreamStackBusLane[22][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane11_strm1_data_valid    ( DownstreamStackBusLane[22][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane12_strm0_ready         ( DownstreamStackBusLane[22][12].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane12_strm0_cntl          ( DownstreamStackBusLane[22][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane12_strm0_data          ( DownstreamStackBusLane[22][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane12_strm0_data_valid    ( DownstreamStackBusLane[22][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane12_strm1_ready         ( DownstreamStackBusLane[22][12].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane12_strm1_cntl          ( DownstreamStackBusLane[22][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane12_strm1_data          ( DownstreamStackBusLane[22][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane12_strm1_data_valid    ( DownstreamStackBusLane[22][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane13_strm0_ready         ( DownstreamStackBusLane[22][13].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane13_strm0_cntl          ( DownstreamStackBusLane[22][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane13_strm0_data          ( DownstreamStackBusLane[22][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane13_strm0_data_valid    ( DownstreamStackBusLane[22][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane13_strm1_ready         ( DownstreamStackBusLane[22][13].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane13_strm1_cntl          ( DownstreamStackBusLane[22][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane13_strm1_data          ( DownstreamStackBusLane[22][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane13_strm1_data_valid    ( DownstreamStackBusLane[22][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane14_strm0_ready         ( DownstreamStackBusLane[22][14].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane14_strm0_cntl          ( DownstreamStackBusLane[22][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane14_strm0_data          ( DownstreamStackBusLane[22][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane14_strm0_data_valid    ( DownstreamStackBusLane[22][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane14_strm1_ready         ( DownstreamStackBusLane[22][14].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane14_strm1_cntl          ( DownstreamStackBusLane[22][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane14_strm1_data          ( DownstreamStackBusLane[22][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane14_strm1_data_valid    ( DownstreamStackBusLane[22][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane15_strm0_ready         ( DownstreamStackBusLane[22][15].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane15_strm0_cntl          ( DownstreamStackBusLane[22][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane15_strm0_data          ( DownstreamStackBusLane[22][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane15_strm0_data_valid    ( DownstreamStackBusLane[22][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane15_strm1_ready         ( DownstreamStackBusLane[22][15].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane15_strm1_cntl          ( DownstreamStackBusLane[22][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane15_strm1_data          ( DownstreamStackBusLane[22][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane15_strm1_data_valid    ( DownstreamStackBusLane[22][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane16_strm0_ready         ( DownstreamStackBusLane[22][16].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane16_strm0_cntl          ( DownstreamStackBusLane[22][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane16_strm0_data          ( DownstreamStackBusLane[22][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane16_strm0_data_valid    ( DownstreamStackBusLane[22][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane16_strm1_ready         ( DownstreamStackBusLane[22][16].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane16_strm1_cntl          ( DownstreamStackBusLane[22][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane16_strm1_data          ( DownstreamStackBusLane[22][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane16_strm1_data_valid    ( DownstreamStackBusLane[22][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane17_strm0_ready         ( DownstreamStackBusLane[22][17].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane17_strm0_cntl          ( DownstreamStackBusLane[22][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane17_strm0_data          ( DownstreamStackBusLane[22][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane17_strm0_data_valid    ( DownstreamStackBusLane[22][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane17_strm1_ready         ( DownstreamStackBusLane[22][17].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane17_strm1_cntl          ( DownstreamStackBusLane[22][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane17_strm1_data          ( DownstreamStackBusLane[22][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane17_strm1_data_valid    ( DownstreamStackBusLane[22][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane18_strm0_ready         ( DownstreamStackBusLane[22][18].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane18_strm0_cntl          ( DownstreamStackBusLane[22][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane18_strm0_data          ( DownstreamStackBusLane[22][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane18_strm0_data_valid    ( DownstreamStackBusLane[22][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane18_strm1_ready         ( DownstreamStackBusLane[22][18].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane18_strm1_cntl          ( DownstreamStackBusLane[22][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane18_strm1_data          ( DownstreamStackBusLane[22][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane18_strm1_data_valid    ( DownstreamStackBusLane[22][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane19_strm0_ready         ( DownstreamStackBusLane[22][19].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane19_strm0_cntl          ( DownstreamStackBusLane[22][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane19_strm0_data          ( DownstreamStackBusLane[22][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane19_strm0_data_valid    ( DownstreamStackBusLane[22][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane19_strm1_ready         ( DownstreamStackBusLane[22][19].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane19_strm1_cntl          ( DownstreamStackBusLane[22][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane19_strm1_data          ( DownstreamStackBusLane[22][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane19_strm1_data_valid    ( DownstreamStackBusLane[22][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane20_strm0_ready         ( DownstreamStackBusLane[22][20].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane20_strm0_cntl          ( DownstreamStackBusLane[22][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane20_strm0_data          ( DownstreamStackBusLane[22][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane20_strm0_data_valid    ( DownstreamStackBusLane[22][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane20_strm1_ready         ( DownstreamStackBusLane[22][20].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane20_strm1_cntl          ( DownstreamStackBusLane[22][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane20_strm1_data          ( DownstreamStackBusLane[22][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane20_strm1_data_valid    ( DownstreamStackBusLane[22][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane21_strm0_ready         ( DownstreamStackBusLane[22][21].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane21_strm0_cntl          ( DownstreamStackBusLane[22][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane21_strm0_data          ( DownstreamStackBusLane[22][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane21_strm0_data_valid    ( DownstreamStackBusLane[22][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane21_strm1_ready         ( DownstreamStackBusLane[22][21].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane21_strm1_cntl          ( DownstreamStackBusLane[22][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane21_strm1_data          ( DownstreamStackBusLane[22][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane21_strm1_data_valid    ( DownstreamStackBusLane[22][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane22_strm0_ready         ( DownstreamStackBusLane[22][22].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane22_strm0_cntl          ( DownstreamStackBusLane[22][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane22_strm0_data          ( DownstreamStackBusLane[22][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane22_strm0_data_valid    ( DownstreamStackBusLane[22][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane22_strm1_ready         ( DownstreamStackBusLane[22][22].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane22_strm1_cntl          ( DownstreamStackBusLane[22][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane22_strm1_data          ( DownstreamStackBusLane[22][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane22_strm1_data_valid    ( DownstreamStackBusLane[22][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane23_strm0_ready         ( DownstreamStackBusLane[22][23].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane23_strm0_cntl          ( DownstreamStackBusLane[22][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane23_strm0_data          ( DownstreamStackBusLane[22][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane23_strm0_data_valid    ( DownstreamStackBusLane[22][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane23_strm1_ready         ( DownstreamStackBusLane[22][23].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane23_strm1_cntl          ( DownstreamStackBusLane[22][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane23_strm1_data          ( DownstreamStackBusLane[22][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane23_strm1_data_valid    ( DownstreamStackBusLane[22][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane24_strm0_ready         ( DownstreamStackBusLane[22][24].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane24_strm0_cntl          ( DownstreamStackBusLane[22][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane24_strm0_data          ( DownstreamStackBusLane[22][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane24_strm0_data_valid    ( DownstreamStackBusLane[22][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane24_strm1_ready         ( DownstreamStackBusLane[22][24].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane24_strm1_cntl          ( DownstreamStackBusLane[22][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane24_strm1_data          ( DownstreamStackBusLane[22][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane24_strm1_data_valid    ( DownstreamStackBusLane[22][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane25_strm0_ready         ( DownstreamStackBusLane[22][25].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane25_strm0_cntl          ( DownstreamStackBusLane[22][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane25_strm0_data          ( DownstreamStackBusLane[22][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane25_strm0_data_valid    ( DownstreamStackBusLane[22][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane25_strm1_ready         ( DownstreamStackBusLane[22][25].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane25_strm1_cntl          ( DownstreamStackBusLane[22][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane25_strm1_data          ( DownstreamStackBusLane[22][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane25_strm1_data_valid    ( DownstreamStackBusLane[22][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane26_strm0_ready         ( DownstreamStackBusLane[22][26].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane26_strm0_cntl          ( DownstreamStackBusLane[22][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane26_strm0_data          ( DownstreamStackBusLane[22][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane26_strm0_data_valid    ( DownstreamStackBusLane[22][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane26_strm1_ready         ( DownstreamStackBusLane[22][26].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane26_strm1_cntl          ( DownstreamStackBusLane[22][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane26_strm1_data          ( DownstreamStackBusLane[22][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane26_strm1_data_valid    ( DownstreamStackBusLane[22][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane27_strm0_ready         ( DownstreamStackBusLane[22][27].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane27_strm0_cntl          ( DownstreamStackBusLane[22][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane27_strm0_data          ( DownstreamStackBusLane[22][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane27_strm0_data_valid    ( DownstreamStackBusLane[22][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane27_strm1_ready         ( DownstreamStackBusLane[22][27].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane27_strm1_cntl          ( DownstreamStackBusLane[22][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane27_strm1_data          ( DownstreamStackBusLane[22][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane27_strm1_data_valid    ( DownstreamStackBusLane[22][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane28_strm0_ready         ( DownstreamStackBusLane[22][28].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane28_strm0_cntl          ( DownstreamStackBusLane[22][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane28_strm0_data          ( DownstreamStackBusLane[22][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane28_strm0_data_valid    ( DownstreamStackBusLane[22][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane28_strm1_ready         ( DownstreamStackBusLane[22][28].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane28_strm1_cntl          ( DownstreamStackBusLane[22][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane28_strm1_data          ( DownstreamStackBusLane[22][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane28_strm1_data_valid    ( DownstreamStackBusLane[22][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane29_strm0_ready         ( DownstreamStackBusLane[22][29].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane29_strm0_cntl          ( DownstreamStackBusLane[22][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane29_strm0_data          ( DownstreamStackBusLane[22][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane29_strm0_data_valid    ( DownstreamStackBusLane[22][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane29_strm1_ready         ( DownstreamStackBusLane[22][29].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane29_strm1_cntl          ( DownstreamStackBusLane[22][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane29_strm1_data          ( DownstreamStackBusLane[22][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane29_strm1_data_valid    ( DownstreamStackBusLane[22][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane30_strm0_ready         ( DownstreamStackBusLane[22][30].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane30_strm0_cntl          ( DownstreamStackBusLane[22][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane30_strm0_data          ( DownstreamStackBusLane[22][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane30_strm0_data_valid    ( DownstreamStackBusLane[22][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane30_strm1_ready         ( DownstreamStackBusLane[22][30].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane30_strm1_cntl          ( DownstreamStackBusLane[22][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane30_strm1_data          ( DownstreamStackBusLane[22][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane30_strm1_data_valid    ( DownstreamStackBusLane[22][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 22, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane31_strm0_ready         ( DownstreamStackBusLane[22][31].pe__std__lane_strm0_ready              ),      
        .std__pe22__lane31_strm0_cntl          ( DownstreamStackBusLane[22][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe22__lane31_strm0_data          ( DownstreamStackBusLane[22][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe22__lane31_strm0_data_valid    ( DownstreamStackBusLane[22][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__std__lane31_strm1_ready         ( DownstreamStackBusLane[22][31].pe__std__lane_strm1_ready              ),      
        .std__pe22__lane31_strm1_cntl          ( DownstreamStackBusLane[22][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe22__lane31_strm1_data          ( DownstreamStackBusLane[22][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe22__lane31_strm1_data_valid    ( DownstreamStackBusLane[22][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane0_strm0_ready         ( DownstreamStackBusLane[23][0].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane0_strm0_cntl          ( DownstreamStackBusLane[23][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane0_strm0_data          ( DownstreamStackBusLane[23][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane0_strm0_data_valid    ( DownstreamStackBusLane[23][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane0_strm1_ready         ( DownstreamStackBusLane[23][0].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane0_strm1_cntl          ( DownstreamStackBusLane[23][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane0_strm1_data          ( DownstreamStackBusLane[23][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane0_strm1_data_valid    ( DownstreamStackBusLane[23][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane1_strm0_ready         ( DownstreamStackBusLane[23][1].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane1_strm0_cntl          ( DownstreamStackBusLane[23][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane1_strm0_data          ( DownstreamStackBusLane[23][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane1_strm0_data_valid    ( DownstreamStackBusLane[23][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane1_strm1_ready         ( DownstreamStackBusLane[23][1].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane1_strm1_cntl          ( DownstreamStackBusLane[23][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane1_strm1_data          ( DownstreamStackBusLane[23][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane1_strm1_data_valid    ( DownstreamStackBusLane[23][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane2_strm0_ready         ( DownstreamStackBusLane[23][2].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane2_strm0_cntl          ( DownstreamStackBusLane[23][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane2_strm0_data          ( DownstreamStackBusLane[23][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane2_strm0_data_valid    ( DownstreamStackBusLane[23][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane2_strm1_ready         ( DownstreamStackBusLane[23][2].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane2_strm1_cntl          ( DownstreamStackBusLane[23][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane2_strm1_data          ( DownstreamStackBusLane[23][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane2_strm1_data_valid    ( DownstreamStackBusLane[23][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane3_strm0_ready         ( DownstreamStackBusLane[23][3].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane3_strm0_cntl          ( DownstreamStackBusLane[23][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane3_strm0_data          ( DownstreamStackBusLane[23][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane3_strm0_data_valid    ( DownstreamStackBusLane[23][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane3_strm1_ready         ( DownstreamStackBusLane[23][3].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane3_strm1_cntl          ( DownstreamStackBusLane[23][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane3_strm1_data          ( DownstreamStackBusLane[23][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane3_strm1_data_valid    ( DownstreamStackBusLane[23][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane4_strm0_ready         ( DownstreamStackBusLane[23][4].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane4_strm0_cntl          ( DownstreamStackBusLane[23][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane4_strm0_data          ( DownstreamStackBusLane[23][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane4_strm0_data_valid    ( DownstreamStackBusLane[23][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane4_strm1_ready         ( DownstreamStackBusLane[23][4].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane4_strm1_cntl          ( DownstreamStackBusLane[23][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane4_strm1_data          ( DownstreamStackBusLane[23][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane4_strm1_data_valid    ( DownstreamStackBusLane[23][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane5_strm0_ready         ( DownstreamStackBusLane[23][5].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane5_strm0_cntl          ( DownstreamStackBusLane[23][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane5_strm0_data          ( DownstreamStackBusLane[23][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane5_strm0_data_valid    ( DownstreamStackBusLane[23][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane5_strm1_ready         ( DownstreamStackBusLane[23][5].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane5_strm1_cntl          ( DownstreamStackBusLane[23][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane5_strm1_data          ( DownstreamStackBusLane[23][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane5_strm1_data_valid    ( DownstreamStackBusLane[23][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane6_strm0_ready         ( DownstreamStackBusLane[23][6].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane6_strm0_cntl          ( DownstreamStackBusLane[23][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane6_strm0_data          ( DownstreamStackBusLane[23][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane6_strm0_data_valid    ( DownstreamStackBusLane[23][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane6_strm1_ready         ( DownstreamStackBusLane[23][6].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane6_strm1_cntl          ( DownstreamStackBusLane[23][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane6_strm1_data          ( DownstreamStackBusLane[23][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane6_strm1_data_valid    ( DownstreamStackBusLane[23][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane7_strm0_ready         ( DownstreamStackBusLane[23][7].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane7_strm0_cntl          ( DownstreamStackBusLane[23][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane7_strm0_data          ( DownstreamStackBusLane[23][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane7_strm0_data_valid    ( DownstreamStackBusLane[23][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane7_strm1_ready         ( DownstreamStackBusLane[23][7].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane7_strm1_cntl          ( DownstreamStackBusLane[23][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane7_strm1_data          ( DownstreamStackBusLane[23][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane7_strm1_data_valid    ( DownstreamStackBusLane[23][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane8_strm0_ready         ( DownstreamStackBusLane[23][8].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane8_strm0_cntl          ( DownstreamStackBusLane[23][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane8_strm0_data          ( DownstreamStackBusLane[23][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane8_strm0_data_valid    ( DownstreamStackBusLane[23][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane8_strm1_ready         ( DownstreamStackBusLane[23][8].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane8_strm1_cntl          ( DownstreamStackBusLane[23][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane8_strm1_data          ( DownstreamStackBusLane[23][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane8_strm1_data_valid    ( DownstreamStackBusLane[23][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane9_strm0_ready         ( DownstreamStackBusLane[23][9].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane9_strm0_cntl          ( DownstreamStackBusLane[23][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane9_strm0_data          ( DownstreamStackBusLane[23][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane9_strm0_data_valid    ( DownstreamStackBusLane[23][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane9_strm1_ready         ( DownstreamStackBusLane[23][9].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane9_strm1_cntl          ( DownstreamStackBusLane[23][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane9_strm1_data          ( DownstreamStackBusLane[23][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane9_strm1_data_valid    ( DownstreamStackBusLane[23][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane10_strm0_ready         ( DownstreamStackBusLane[23][10].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane10_strm0_cntl          ( DownstreamStackBusLane[23][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane10_strm0_data          ( DownstreamStackBusLane[23][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane10_strm0_data_valid    ( DownstreamStackBusLane[23][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane10_strm1_ready         ( DownstreamStackBusLane[23][10].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane10_strm1_cntl          ( DownstreamStackBusLane[23][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane10_strm1_data          ( DownstreamStackBusLane[23][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane10_strm1_data_valid    ( DownstreamStackBusLane[23][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane11_strm0_ready         ( DownstreamStackBusLane[23][11].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane11_strm0_cntl          ( DownstreamStackBusLane[23][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane11_strm0_data          ( DownstreamStackBusLane[23][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane11_strm0_data_valid    ( DownstreamStackBusLane[23][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane11_strm1_ready         ( DownstreamStackBusLane[23][11].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane11_strm1_cntl          ( DownstreamStackBusLane[23][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane11_strm1_data          ( DownstreamStackBusLane[23][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane11_strm1_data_valid    ( DownstreamStackBusLane[23][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane12_strm0_ready         ( DownstreamStackBusLane[23][12].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane12_strm0_cntl          ( DownstreamStackBusLane[23][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane12_strm0_data          ( DownstreamStackBusLane[23][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane12_strm0_data_valid    ( DownstreamStackBusLane[23][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane12_strm1_ready         ( DownstreamStackBusLane[23][12].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane12_strm1_cntl          ( DownstreamStackBusLane[23][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane12_strm1_data          ( DownstreamStackBusLane[23][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane12_strm1_data_valid    ( DownstreamStackBusLane[23][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane13_strm0_ready         ( DownstreamStackBusLane[23][13].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane13_strm0_cntl          ( DownstreamStackBusLane[23][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane13_strm0_data          ( DownstreamStackBusLane[23][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane13_strm0_data_valid    ( DownstreamStackBusLane[23][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane13_strm1_ready         ( DownstreamStackBusLane[23][13].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane13_strm1_cntl          ( DownstreamStackBusLane[23][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane13_strm1_data          ( DownstreamStackBusLane[23][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane13_strm1_data_valid    ( DownstreamStackBusLane[23][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane14_strm0_ready         ( DownstreamStackBusLane[23][14].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane14_strm0_cntl          ( DownstreamStackBusLane[23][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane14_strm0_data          ( DownstreamStackBusLane[23][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane14_strm0_data_valid    ( DownstreamStackBusLane[23][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane14_strm1_ready         ( DownstreamStackBusLane[23][14].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane14_strm1_cntl          ( DownstreamStackBusLane[23][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane14_strm1_data          ( DownstreamStackBusLane[23][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane14_strm1_data_valid    ( DownstreamStackBusLane[23][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane15_strm0_ready         ( DownstreamStackBusLane[23][15].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane15_strm0_cntl          ( DownstreamStackBusLane[23][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane15_strm0_data          ( DownstreamStackBusLane[23][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane15_strm0_data_valid    ( DownstreamStackBusLane[23][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane15_strm1_ready         ( DownstreamStackBusLane[23][15].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane15_strm1_cntl          ( DownstreamStackBusLane[23][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane15_strm1_data          ( DownstreamStackBusLane[23][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane15_strm1_data_valid    ( DownstreamStackBusLane[23][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane16_strm0_ready         ( DownstreamStackBusLane[23][16].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane16_strm0_cntl          ( DownstreamStackBusLane[23][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane16_strm0_data          ( DownstreamStackBusLane[23][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane16_strm0_data_valid    ( DownstreamStackBusLane[23][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane16_strm1_ready         ( DownstreamStackBusLane[23][16].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane16_strm1_cntl          ( DownstreamStackBusLane[23][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane16_strm1_data          ( DownstreamStackBusLane[23][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane16_strm1_data_valid    ( DownstreamStackBusLane[23][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane17_strm0_ready         ( DownstreamStackBusLane[23][17].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane17_strm0_cntl          ( DownstreamStackBusLane[23][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane17_strm0_data          ( DownstreamStackBusLane[23][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane17_strm0_data_valid    ( DownstreamStackBusLane[23][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane17_strm1_ready         ( DownstreamStackBusLane[23][17].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane17_strm1_cntl          ( DownstreamStackBusLane[23][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane17_strm1_data          ( DownstreamStackBusLane[23][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane17_strm1_data_valid    ( DownstreamStackBusLane[23][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane18_strm0_ready         ( DownstreamStackBusLane[23][18].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane18_strm0_cntl          ( DownstreamStackBusLane[23][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane18_strm0_data          ( DownstreamStackBusLane[23][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane18_strm0_data_valid    ( DownstreamStackBusLane[23][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane18_strm1_ready         ( DownstreamStackBusLane[23][18].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane18_strm1_cntl          ( DownstreamStackBusLane[23][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane18_strm1_data          ( DownstreamStackBusLane[23][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane18_strm1_data_valid    ( DownstreamStackBusLane[23][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane19_strm0_ready         ( DownstreamStackBusLane[23][19].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane19_strm0_cntl          ( DownstreamStackBusLane[23][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane19_strm0_data          ( DownstreamStackBusLane[23][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane19_strm0_data_valid    ( DownstreamStackBusLane[23][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane19_strm1_ready         ( DownstreamStackBusLane[23][19].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane19_strm1_cntl          ( DownstreamStackBusLane[23][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane19_strm1_data          ( DownstreamStackBusLane[23][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane19_strm1_data_valid    ( DownstreamStackBusLane[23][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane20_strm0_ready         ( DownstreamStackBusLane[23][20].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane20_strm0_cntl          ( DownstreamStackBusLane[23][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane20_strm0_data          ( DownstreamStackBusLane[23][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane20_strm0_data_valid    ( DownstreamStackBusLane[23][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane20_strm1_ready         ( DownstreamStackBusLane[23][20].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane20_strm1_cntl          ( DownstreamStackBusLane[23][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane20_strm1_data          ( DownstreamStackBusLane[23][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane20_strm1_data_valid    ( DownstreamStackBusLane[23][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane21_strm0_ready         ( DownstreamStackBusLane[23][21].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane21_strm0_cntl          ( DownstreamStackBusLane[23][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane21_strm0_data          ( DownstreamStackBusLane[23][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane21_strm0_data_valid    ( DownstreamStackBusLane[23][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane21_strm1_ready         ( DownstreamStackBusLane[23][21].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane21_strm1_cntl          ( DownstreamStackBusLane[23][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane21_strm1_data          ( DownstreamStackBusLane[23][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane21_strm1_data_valid    ( DownstreamStackBusLane[23][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane22_strm0_ready         ( DownstreamStackBusLane[23][22].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane22_strm0_cntl          ( DownstreamStackBusLane[23][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane22_strm0_data          ( DownstreamStackBusLane[23][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane22_strm0_data_valid    ( DownstreamStackBusLane[23][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane22_strm1_ready         ( DownstreamStackBusLane[23][22].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane22_strm1_cntl          ( DownstreamStackBusLane[23][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane22_strm1_data          ( DownstreamStackBusLane[23][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane22_strm1_data_valid    ( DownstreamStackBusLane[23][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane23_strm0_ready         ( DownstreamStackBusLane[23][23].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane23_strm0_cntl          ( DownstreamStackBusLane[23][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane23_strm0_data          ( DownstreamStackBusLane[23][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane23_strm0_data_valid    ( DownstreamStackBusLane[23][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane23_strm1_ready         ( DownstreamStackBusLane[23][23].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane23_strm1_cntl          ( DownstreamStackBusLane[23][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane23_strm1_data          ( DownstreamStackBusLane[23][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane23_strm1_data_valid    ( DownstreamStackBusLane[23][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane24_strm0_ready         ( DownstreamStackBusLane[23][24].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane24_strm0_cntl          ( DownstreamStackBusLane[23][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane24_strm0_data          ( DownstreamStackBusLane[23][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane24_strm0_data_valid    ( DownstreamStackBusLane[23][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane24_strm1_ready         ( DownstreamStackBusLane[23][24].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane24_strm1_cntl          ( DownstreamStackBusLane[23][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane24_strm1_data          ( DownstreamStackBusLane[23][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane24_strm1_data_valid    ( DownstreamStackBusLane[23][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane25_strm0_ready         ( DownstreamStackBusLane[23][25].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane25_strm0_cntl          ( DownstreamStackBusLane[23][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane25_strm0_data          ( DownstreamStackBusLane[23][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane25_strm0_data_valid    ( DownstreamStackBusLane[23][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane25_strm1_ready         ( DownstreamStackBusLane[23][25].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane25_strm1_cntl          ( DownstreamStackBusLane[23][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane25_strm1_data          ( DownstreamStackBusLane[23][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane25_strm1_data_valid    ( DownstreamStackBusLane[23][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane26_strm0_ready         ( DownstreamStackBusLane[23][26].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane26_strm0_cntl          ( DownstreamStackBusLane[23][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane26_strm0_data          ( DownstreamStackBusLane[23][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane26_strm0_data_valid    ( DownstreamStackBusLane[23][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane26_strm1_ready         ( DownstreamStackBusLane[23][26].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane26_strm1_cntl          ( DownstreamStackBusLane[23][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane26_strm1_data          ( DownstreamStackBusLane[23][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane26_strm1_data_valid    ( DownstreamStackBusLane[23][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane27_strm0_ready         ( DownstreamStackBusLane[23][27].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane27_strm0_cntl          ( DownstreamStackBusLane[23][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane27_strm0_data          ( DownstreamStackBusLane[23][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane27_strm0_data_valid    ( DownstreamStackBusLane[23][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane27_strm1_ready         ( DownstreamStackBusLane[23][27].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane27_strm1_cntl          ( DownstreamStackBusLane[23][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane27_strm1_data          ( DownstreamStackBusLane[23][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane27_strm1_data_valid    ( DownstreamStackBusLane[23][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane28_strm0_ready         ( DownstreamStackBusLane[23][28].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane28_strm0_cntl          ( DownstreamStackBusLane[23][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane28_strm0_data          ( DownstreamStackBusLane[23][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane28_strm0_data_valid    ( DownstreamStackBusLane[23][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane28_strm1_ready         ( DownstreamStackBusLane[23][28].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane28_strm1_cntl          ( DownstreamStackBusLane[23][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane28_strm1_data          ( DownstreamStackBusLane[23][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane28_strm1_data_valid    ( DownstreamStackBusLane[23][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane29_strm0_ready         ( DownstreamStackBusLane[23][29].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane29_strm0_cntl          ( DownstreamStackBusLane[23][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane29_strm0_data          ( DownstreamStackBusLane[23][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane29_strm0_data_valid    ( DownstreamStackBusLane[23][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane29_strm1_ready         ( DownstreamStackBusLane[23][29].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane29_strm1_cntl          ( DownstreamStackBusLane[23][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane29_strm1_data          ( DownstreamStackBusLane[23][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane29_strm1_data_valid    ( DownstreamStackBusLane[23][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane30_strm0_ready         ( DownstreamStackBusLane[23][30].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane30_strm0_cntl          ( DownstreamStackBusLane[23][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane30_strm0_data          ( DownstreamStackBusLane[23][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane30_strm0_data_valid    ( DownstreamStackBusLane[23][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane30_strm1_ready         ( DownstreamStackBusLane[23][30].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane30_strm1_cntl          ( DownstreamStackBusLane[23][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane30_strm1_data          ( DownstreamStackBusLane[23][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane30_strm1_data_valid    ( DownstreamStackBusLane[23][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 23, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane31_strm0_ready         ( DownstreamStackBusLane[23][31].pe__std__lane_strm0_ready              ),      
        .std__pe23__lane31_strm0_cntl          ( DownstreamStackBusLane[23][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe23__lane31_strm0_data          ( DownstreamStackBusLane[23][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe23__lane31_strm0_data_valid    ( DownstreamStackBusLane[23][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__std__lane31_strm1_ready         ( DownstreamStackBusLane[23][31].pe__std__lane_strm1_ready              ),      
        .std__pe23__lane31_strm1_cntl          ( DownstreamStackBusLane[23][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe23__lane31_strm1_data          ( DownstreamStackBusLane[23][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe23__lane31_strm1_data_valid    ( DownstreamStackBusLane[23][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane0_strm0_ready         ( DownstreamStackBusLane[24][0].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane0_strm0_cntl          ( DownstreamStackBusLane[24][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane0_strm0_data          ( DownstreamStackBusLane[24][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane0_strm0_data_valid    ( DownstreamStackBusLane[24][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane0_strm1_ready         ( DownstreamStackBusLane[24][0].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane0_strm1_cntl          ( DownstreamStackBusLane[24][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane0_strm1_data          ( DownstreamStackBusLane[24][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane0_strm1_data_valid    ( DownstreamStackBusLane[24][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane1_strm0_ready         ( DownstreamStackBusLane[24][1].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane1_strm0_cntl          ( DownstreamStackBusLane[24][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane1_strm0_data          ( DownstreamStackBusLane[24][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane1_strm0_data_valid    ( DownstreamStackBusLane[24][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane1_strm1_ready         ( DownstreamStackBusLane[24][1].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane1_strm1_cntl          ( DownstreamStackBusLane[24][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane1_strm1_data          ( DownstreamStackBusLane[24][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane1_strm1_data_valid    ( DownstreamStackBusLane[24][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane2_strm0_ready         ( DownstreamStackBusLane[24][2].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane2_strm0_cntl          ( DownstreamStackBusLane[24][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane2_strm0_data          ( DownstreamStackBusLane[24][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane2_strm0_data_valid    ( DownstreamStackBusLane[24][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane2_strm1_ready         ( DownstreamStackBusLane[24][2].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane2_strm1_cntl          ( DownstreamStackBusLane[24][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane2_strm1_data          ( DownstreamStackBusLane[24][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane2_strm1_data_valid    ( DownstreamStackBusLane[24][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane3_strm0_ready         ( DownstreamStackBusLane[24][3].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane3_strm0_cntl          ( DownstreamStackBusLane[24][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane3_strm0_data          ( DownstreamStackBusLane[24][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane3_strm0_data_valid    ( DownstreamStackBusLane[24][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane3_strm1_ready         ( DownstreamStackBusLane[24][3].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane3_strm1_cntl          ( DownstreamStackBusLane[24][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane3_strm1_data          ( DownstreamStackBusLane[24][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane3_strm1_data_valid    ( DownstreamStackBusLane[24][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane4_strm0_ready         ( DownstreamStackBusLane[24][4].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane4_strm0_cntl          ( DownstreamStackBusLane[24][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane4_strm0_data          ( DownstreamStackBusLane[24][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane4_strm0_data_valid    ( DownstreamStackBusLane[24][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane4_strm1_ready         ( DownstreamStackBusLane[24][4].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane4_strm1_cntl          ( DownstreamStackBusLane[24][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane4_strm1_data          ( DownstreamStackBusLane[24][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane4_strm1_data_valid    ( DownstreamStackBusLane[24][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane5_strm0_ready         ( DownstreamStackBusLane[24][5].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane5_strm0_cntl          ( DownstreamStackBusLane[24][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane5_strm0_data          ( DownstreamStackBusLane[24][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane5_strm0_data_valid    ( DownstreamStackBusLane[24][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane5_strm1_ready         ( DownstreamStackBusLane[24][5].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane5_strm1_cntl          ( DownstreamStackBusLane[24][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane5_strm1_data          ( DownstreamStackBusLane[24][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane5_strm1_data_valid    ( DownstreamStackBusLane[24][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane6_strm0_ready         ( DownstreamStackBusLane[24][6].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane6_strm0_cntl          ( DownstreamStackBusLane[24][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane6_strm0_data          ( DownstreamStackBusLane[24][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane6_strm0_data_valid    ( DownstreamStackBusLane[24][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane6_strm1_ready         ( DownstreamStackBusLane[24][6].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane6_strm1_cntl          ( DownstreamStackBusLane[24][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane6_strm1_data          ( DownstreamStackBusLane[24][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane6_strm1_data_valid    ( DownstreamStackBusLane[24][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane7_strm0_ready         ( DownstreamStackBusLane[24][7].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane7_strm0_cntl          ( DownstreamStackBusLane[24][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane7_strm0_data          ( DownstreamStackBusLane[24][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane7_strm0_data_valid    ( DownstreamStackBusLane[24][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane7_strm1_ready         ( DownstreamStackBusLane[24][7].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane7_strm1_cntl          ( DownstreamStackBusLane[24][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane7_strm1_data          ( DownstreamStackBusLane[24][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane7_strm1_data_valid    ( DownstreamStackBusLane[24][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane8_strm0_ready         ( DownstreamStackBusLane[24][8].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane8_strm0_cntl          ( DownstreamStackBusLane[24][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane8_strm0_data          ( DownstreamStackBusLane[24][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane8_strm0_data_valid    ( DownstreamStackBusLane[24][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane8_strm1_ready         ( DownstreamStackBusLane[24][8].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane8_strm1_cntl          ( DownstreamStackBusLane[24][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane8_strm1_data          ( DownstreamStackBusLane[24][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane8_strm1_data_valid    ( DownstreamStackBusLane[24][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane9_strm0_ready         ( DownstreamStackBusLane[24][9].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane9_strm0_cntl          ( DownstreamStackBusLane[24][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane9_strm0_data          ( DownstreamStackBusLane[24][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane9_strm0_data_valid    ( DownstreamStackBusLane[24][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane9_strm1_ready         ( DownstreamStackBusLane[24][9].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane9_strm1_cntl          ( DownstreamStackBusLane[24][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane9_strm1_data          ( DownstreamStackBusLane[24][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane9_strm1_data_valid    ( DownstreamStackBusLane[24][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane10_strm0_ready         ( DownstreamStackBusLane[24][10].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane10_strm0_cntl          ( DownstreamStackBusLane[24][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane10_strm0_data          ( DownstreamStackBusLane[24][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane10_strm0_data_valid    ( DownstreamStackBusLane[24][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane10_strm1_ready         ( DownstreamStackBusLane[24][10].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane10_strm1_cntl          ( DownstreamStackBusLane[24][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane10_strm1_data          ( DownstreamStackBusLane[24][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane10_strm1_data_valid    ( DownstreamStackBusLane[24][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane11_strm0_ready         ( DownstreamStackBusLane[24][11].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane11_strm0_cntl          ( DownstreamStackBusLane[24][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane11_strm0_data          ( DownstreamStackBusLane[24][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane11_strm0_data_valid    ( DownstreamStackBusLane[24][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane11_strm1_ready         ( DownstreamStackBusLane[24][11].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane11_strm1_cntl          ( DownstreamStackBusLane[24][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane11_strm1_data          ( DownstreamStackBusLane[24][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane11_strm1_data_valid    ( DownstreamStackBusLane[24][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane12_strm0_ready         ( DownstreamStackBusLane[24][12].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane12_strm0_cntl          ( DownstreamStackBusLane[24][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane12_strm0_data          ( DownstreamStackBusLane[24][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane12_strm0_data_valid    ( DownstreamStackBusLane[24][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane12_strm1_ready         ( DownstreamStackBusLane[24][12].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane12_strm1_cntl          ( DownstreamStackBusLane[24][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane12_strm1_data          ( DownstreamStackBusLane[24][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane12_strm1_data_valid    ( DownstreamStackBusLane[24][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane13_strm0_ready         ( DownstreamStackBusLane[24][13].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane13_strm0_cntl          ( DownstreamStackBusLane[24][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane13_strm0_data          ( DownstreamStackBusLane[24][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane13_strm0_data_valid    ( DownstreamStackBusLane[24][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane13_strm1_ready         ( DownstreamStackBusLane[24][13].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane13_strm1_cntl          ( DownstreamStackBusLane[24][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane13_strm1_data          ( DownstreamStackBusLane[24][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane13_strm1_data_valid    ( DownstreamStackBusLane[24][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane14_strm0_ready         ( DownstreamStackBusLane[24][14].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane14_strm0_cntl          ( DownstreamStackBusLane[24][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane14_strm0_data          ( DownstreamStackBusLane[24][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane14_strm0_data_valid    ( DownstreamStackBusLane[24][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane14_strm1_ready         ( DownstreamStackBusLane[24][14].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane14_strm1_cntl          ( DownstreamStackBusLane[24][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane14_strm1_data          ( DownstreamStackBusLane[24][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane14_strm1_data_valid    ( DownstreamStackBusLane[24][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane15_strm0_ready         ( DownstreamStackBusLane[24][15].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane15_strm0_cntl          ( DownstreamStackBusLane[24][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane15_strm0_data          ( DownstreamStackBusLane[24][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane15_strm0_data_valid    ( DownstreamStackBusLane[24][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane15_strm1_ready         ( DownstreamStackBusLane[24][15].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane15_strm1_cntl          ( DownstreamStackBusLane[24][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane15_strm1_data          ( DownstreamStackBusLane[24][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane15_strm1_data_valid    ( DownstreamStackBusLane[24][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane16_strm0_ready         ( DownstreamStackBusLane[24][16].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane16_strm0_cntl          ( DownstreamStackBusLane[24][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane16_strm0_data          ( DownstreamStackBusLane[24][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane16_strm0_data_valid    ( DownstreamStackBusLane[24][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane16_strm1_ready         ( DownstreamStackBusLane[24][16].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane16_strm1_cntl          ( DownstreamStackBusLane[24][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane16_strm1_data          ( DownstreamStackBusLane[24][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane16_strm1_data_valid    ( DownstreamStackBusLane[24][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane17_strm0_ready         ( DownstreamStackBusLane[24][17].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane17_strm0_cntl          ( DownstreamStackBusLane[24][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane17_strm0_data          ( DownstreamStackBusLane[24][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane17_strm0_data_valid    ( DownstreamStackBusLane[24][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane17_strm1_ready         ( DownstreamStackBusLane[24][17].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane17_strm1_cntl          ( DownstreamStackBusLane[24][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane17_strm1_data          ( DownstreamStackBusLane[24][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane17_strm1_data_valid    ( DownstreamStackBusLane[24][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane18_strm0_ready         ( DownstreamStackBusLane[24][18].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane18_strm0_cntl          ( DownstreamStackBusLane[24][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane18_strm0_data          ( DownstreamStackBusLane[24][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane18_strm0_data_valid    ( DownstreamStackBusLane[24][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane18_strm1_ready         ( DownstreamStackBusLane[24][18].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane18_strm1_cntl          ( DownstreamStackBusLane[24][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane18_strm1_data          ( DownstreamStackBusLane[24][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane18_strm1_data_valid    ( DownstreamStackBusLane[24][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane19_strm0_ready         ( DownstreamStackBusLane[24][19].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane19_strm0_cntl          ( DownstreamStackBusLane[24][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane19_strm0_data          ( DownstreamStackBusLane[24][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane19_strm0_data_valid    ( DownstreamStackBusLane[24][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane19_strm1_ready         ( DownstreamStackBusLane[24][19].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane19_strm1_cntl          ( DownstreamStackBusLane[24][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane19_strm1_data          ( DownstreamStackBusLane[24][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane19_strm1_data_valid    ( DownstreamStackBusLane[24][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane20_strm0_ready         ( DownstreamStackBusLane[24][20].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane20_strm0_cntl          ( DownstreamStackBusLane[24][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane20_strm0_data          ( DownstreamStackBusLane[24][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane20_strm0_data_valid    ( DownstreamStackBusLane[24][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane20_strm1_ready         ( DownstreamStackBusLane[24][20].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane20_strm1_cntl          ( DownstreamStackBusLane[24][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane20_strm1_data          ( DownstreamStackBusLane[24][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane20_strm1_data_valid    ( DownstreamStackBusLane[24][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane21_strm0_ready         ( DownstreamStackBusLane[24][21].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane21_strm0_cntl          ( DownstreamStackBusLane[24][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane21_strm0_data          ( DownstreamStackBusLane[24][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane21_strm0_data_valid    ( DownstreamStackBusLane[24][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane21_strm1_ready         ( DownstreamStackBusLane[24][21].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane21_strm1_cntl          ( DownstreamStackBusLane[24][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane21_strm1_data          ( DownstreamStackBusLane[24][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane21_strm1_data_valid    ( DownstreamStackBusLane[24][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane22_strm0_ready         ( DownstreamStackBusLane[24][22].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane22_strm0_cntl          ( DownstreamStackBusLane[24][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane22_strm0_data          ( DownstreamStackBusLane[24][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane22_strm0_data_valid    ( DownstreamStackBusLane[24][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane22_strm1_ready         ( DownstreamStackBusLane[24][22].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane22_strm1_cntl          ( DownstreamStackBusLane[24][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane22_strm1_data          ( DownstreamStackBusLane[24][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane22_strm1_data_valid    ( DownstreamStackBusLane[24][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane23_strm0_ready         ( DownstreamStackBusLane[24][23].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane23_strm0_cntl          ( DownstreamStackBusLane[24][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane23_strm0_data          ( DownstreamStackBusLane[24][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane23_strm0_data_valid    ( DownstreamStackBusLane[24][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane23_strm1_ready         ( DownstreamStackBusLane[24][23].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane23_strm1_cntl          ( DownstreamStackBusLane[24][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane23_strm1_data          ( DownstreamStackBusLane[24][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane23_strm1_data_valid    ( DownstreamStackBusLane[24][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane24_strm0_ready         ( DownstreamStackBusLane[24][24].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane24_strm0_cntl          ( DownstreamStackBusLane[24][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane24_strm0_data          ( DownstreamStackBusLane[24][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane24_strm0_data_valid    ( DownstreamStackBusLane[24][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane24_strm1_ready         ( DownstreamStackBusLane[24][24].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane24_strm1_cntl          ( DownstreamStackBusLane[24][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane24_strm1_data          ( DownstreamStackBusLane[24][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane24_strm1_data_valid    ( DownstreamStackBusLane[24][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane25_strm0_ready         ( DownstreamStackBusLane[24][25].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane25_strm0_cntl          ( DownstreamStackBusLane[24][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane25_strm0_data          ( DownstreamStackBusLane[24][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane25_strm0_data_valid    ( DownstreamStackBusLane[24][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane25_strm1_ready         ( DownstreamStackBusLane[24][25].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane25_strm1_cntl          ( DownstreamStackBusLane[24][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane25_strm1_data          ( DownstreamStackBusLane[24][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane25_strm1_data_valid    ( DownstreamStackBusLane[24][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane26_strm0_ready         ( DownstreamStackBusLane[24][26].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane26_strm0_cntl          ( DownstreamStackBusLane[24][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane26_strm0_data          ( DownstreamStackBusLane[24][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane26_strm0_data_valid    ( DownstreamStackBusLane[24][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane26_strm1_ready         ( DownstreamStackBusLane[24][26].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane26_strm1_cntl          ( DownstreamStackBusLane[24][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane26_strm1_data          ( DownstreamStackBusLane[24][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane26_strm1_data_valid    ( DownstreamStackBusLane[24][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane27_strm0_ready         ( DownstreamStackBusLane[24][27].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane27_strm0_cntl          ( DownstreamStackBusLane[24][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane27_strm0_data          ( DownstreamStackBusLane[24][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane27_strm0_data_valid    ( DownstreamStackBusLane[24][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane27_strm1_ready         ( DownstreamStackBusLane[24][27].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane27_strm1_cntl          ( DownstreamStackBusLane[24][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane27_strm1_data          ( DownstreamStackBusLane[24][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane27_strm1_data_valid    ( DownstreamStackBusLane[24][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane28_strm0_ready         ( DownstreamStackBusLane[24][28].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane28_strm0_cntl          ( DownstreamStackBusLane[24][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane28_strm0_data          ( DownstreamStackBusLane[24][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane28_strm0_data_valid    ( DownstreamStackBusLane[24][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane28_strm1_ready         ( DownstreamStackBusLane[24][28].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane28_strm1_cntl          ( DownstreamStackBusLane[24][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane28_strm1_data          ( DownstreamStackBusLane[24][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane28_strm1_data_valid    ( DownstreamStackBusLane[24][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane29_strm0_ready         ( DownstreamStackBusLane[24][29].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane29_strm0_cntl          ( DownstreamStackBusLane[24][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane29_strm0_data          ( DownstreamStackBusLane[24][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane29_strm0_data_valid    ( DownstreamStackBusLane[24][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane29_strm1_ready         ( DownstreamStackBusLane[24][29].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane29_strm1_cntl          ( DownstreamStackBusLane[24][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane29_strm1_data          ( DownstreamStackBusLane[24][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane29_strm1_data_valid    ( DownstreamStackBusLane[24][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane30_strm0_ready         ( DownstreamStackBusLane[24][30].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane30_strm0_cntl          ( DownstreamStackBusLane[24][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane30_strm0_data          ( DownstreamStackBusLane[24][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane30_strm0_data_valid    ( DownstreamStackBusLane[24][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane30_strm1_ready         ( DownstreamStackBusLane[24][30].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane30_strm1_cntl          ( DownstreamStackBusLane[24][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane30_strm1_data          ( DownstreamStackBusLane[24][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane30_strm1_data_valid    ( DownstreamStackBusLane[24][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 24, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane31_strm0_ready         ( DownstreamStackBusLane[24][31].pe__std__lane_strm0_ready              ),      
        .std__pe24__lane31_strm0_cntl          ( DownstreamStackBusLane[24][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe24__lane31_strm0_data          ( DownstreamStackBusLane[24][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe24__lane31_strm0_data_valid    ( DownstreamStackBusLane[24][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__std__lane31_strm1_ready         ( DownstreamStackBusLane[24][31].pe__std__lane_strm1_ready              ),      
        .std__pe24__lane31_strm1_cntl          ( DownstreamStackBusLane[24][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe24__lane31_strm1_data          ( DownstreamStackBusLane[24][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe24__lane31_strm1_data_valid    ( DownstreamStackBusLane[24][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane0_strm0_ready         ( DownstreamStackBusLane[25][0].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane0_strm0_cntl          ( DownstreamStackBusLane[25][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane0_strm0_data          ( DownstreamStackBusLane[25][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane0_strm0_data_valid    ( DownstreamStackBusLane[25][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane0_strm1_ready         ( DownstreamStackBusLane[25][0].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane0_strm1_cntl          ( DownstreamStackBusLane[25][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane0_strm1_data          ( DownstreamStackBusLane[25][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane0_strm1_data_valid    ( DownstreamStackBusLane[25][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane1_strm0_ready         ( DownstreamStackBusLane[25][1].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane1_strm0_cntl          ( DownstreamStackBusLane[25][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane1_strm0_data          ( DownstreamStackBusLane[25][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane1_strm0_data_valid    ( DownstreamStackBusLane[25][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane1_strm1_ready         ( DownstreamStackBusLane[25][1].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane1_strm1_cntl          ( DownstreamStackBusLane[25][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane1_strm1_data          ( DownstreamStackBusLane[25][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane1_strm1_data_valid    ( DownstreamStackBusLane[25][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane2_strm0_ready         ( DownstreamStackBusLane[25][2].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane2_strm0_cntl          ( DownstreamStackBusLane[25][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane2_strm0_data          ( DownstreamStackBusLane[25][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane2_strm0_data_valid    ( DownstreamStackBusLane[25][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane2_strm1_ready         ( DownstreamStackBusLane[25][2].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane2_strm1_cntl          ( DownstreamStackBusLane[25][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane2_strm1_data          ( DownstreamStackBusLane[25][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane2_strm1_data_valid    ( DownstreamStackBusLane[25][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane3_strm0_ready         ( DownstreamStackBusLane[25][3].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane3_strm0_cntl          ( DownstreamStackBusLane[25][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane3_strm0_data          ( DownstreamStackBusLane[25][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane3_strm0_data_valid    ( DownstreamStackBusLane[25][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane3_strm1_ready         ( DownstreamStackBusLane[25][3].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane3_strm1_cntl          ( DownstreamStackBusLane[25][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane3_strm1_data          ( DownstreamStackBusLane[25][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane3_strm1_data_valid    ( DownstreamStackBusLane[25][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane4_strm0_ready         ( DownstreamStackBusLane[25][4].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane4_strm0_cntl          ( DownstreamStackBusLane[25][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane4_strm0_data          ( DownstreamStackBusLane[25][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane4_strm0_data_valid    ( DownstreamStackBusLane[25][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane4_strm1_ready         ( DownstreamStackBusLane[25][4].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane4_strm1_cntl          ( DownstreamStackBusLane[25][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane4_strm1_data          ( DownstreamStackBusLane[25][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane4_strm1_data_valid    ( DownstreamStackBusLane[25][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane5_strm0_ready         ( DownstreamStackBusLane[25][5].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane5_strm0_cntl          ( DownstreamStackBusLane[25][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane5_strm0_data          ( DownstreamStackBusLane[25][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane5_strm0_data_valid    ( DownstreamStackBusLane[25][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane5_strm1_ready         ( DownstreamStackBusLane[25][5].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane5_strm1_cntl          ( DownstreamStackBusLane[25][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane5_strm1_data          ( DownstreamStackBusLane[25][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane5_strm1_data_valid    ( DownstreamStackBusLane[25][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane6_strm0_ready         ( DownstreamStackBusLane[25][6].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane6_strm0_cntl          ( DownstreamStackBusLane[25][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane6_strm0_data          ( DownstreamStackBusLane[25][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane6_strm0_data_valid    ( DownstreamStackBusLane[25][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane6_strm1_ready         ( DownstreamStackBusLane[25][6].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane6_strm1_cntl          ( DownstreamStackBusLane[25][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane6_strm1_data          ( DownstreamStackBusLane[25][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane6_strm1_data_valid    ( DownstreamStackBusLane[25][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane7_strm0_ready         ( DownstreamStackBusLane[25][7].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane7_strm0_cntl          ( DownstreamStackBusLane[25][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane7_strm0_data          ( DownstreamStackBusLane[25][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane7_strm0_data_valid    ( DownstreamStackBusLane[25][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane7_strm1_ready         ( DownstreamStackBusLane[25][7].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane7_strm1_cntl          ( DownstreamStackBusLane[25][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane7_strm1_data          ( DownstreamStackBusLane[25][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane7_strm1_data_valid    ( DownstreamStackBusLane[25][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane8_strm0_ready         ( DownstreamStackBusLane[25][8].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane8_strm0_cntl          ( DownstreamStackBusLane[25][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane8_strm0_data          ( DownstreamStackBusLane[25][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane8_strm0_data_valid    ( DownstreamStackBusLane[25][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane8_strm1_ready         ( DownstreamStackBusLane[25][8].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane8_strm1_cntl          ( DownstreamStackBusLane[25][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane8_strm1_data          ( DownstreamStackBusLane[25][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane8_strm1_data_valid    ( DownstreamStackBusLane[25][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane9_strm0_ready         ( DownstreamStackBusLane[25][9].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane9_strm0_cntl          ( DownstreamStackBusLane[25][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane9_strm0_data          ( DownstreamStackBusLane[25][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane9_strm0_data_valid    ( DownstreamStackBusLane[25][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane9_strm1_ready         ( DownstreamStackBusLane[25][9].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane9_strm1_cntl          ( DownstreamStackBusLane[25][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane9_strm1_data          ( DownstreamStackBusLane[25][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane9_strm1_data_valid    ( DownstreamStackBusLane[25][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane10_strm0_ready         ( DownstreamStackBusLane[25][10].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane10_strm0_cntl          ( DownstreamStackBusLane[25][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane10_strm0_data          ( DownstreamStackBusLane[25][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane10_strm0_data_valid    ( DownstreamStackBusLane[25][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane10_strm1_ready         ( DownstreamStackBusLane[25][10].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane10_strm1_cntl          ( DownstreamStackBusLane[25][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane10_strm1_data          ( DownstreamStackBusLane[25][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane10_strm1_data_valid    ( DownstreamStackBusLane[25][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane11_strm0_ready         ( DownstreamStackBusLane[25][11].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane11_strm0_cntl          ( DownstreamStackBusLane[25][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane11_strm0_data          ( DownstreamStackBusLane[25][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane11_strm0_data_valid    ( DownstreamStackBusLane[25][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane11_strm1_ready         ( DownstreamStackBusLane[25][11].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane11_strm1_cntl          ( DownstreamStackBusLane[25][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane11_strm1_data          ( DownstreamStackBusLane[25][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane11_strm1_data_valid    ( DownstreamStackBusLane[25][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane12_strm0_ready         ( DownstreamStackBusLane[25][12].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane12_strm0_cntl          ( DownstreamStackBusLane[25][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane12_strm0_data          ( DownstreamStackBusLane[25][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane12_strm0_data_valid    ( DownstreamStackBusLane[25][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane12_strm1_ready         ( DownstreamStackBusLane[25][12].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane12_strm1_cntl          ( DownstreamStackBusLane[25][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane12_strm1_data          ( DownstreamStackBusLane[25][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane12_strm1_data_valid    ( DownstreamStackBusLane[25][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane13_strm0_ready         ( DownstreamStackBusLane[25][13].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane13_strm0_cntl          ( DownstreamStackBusLane[25][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane13_strm0_data          ( DownstreamStackBusLane[25][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane13_strm0_data_valid    ( DownstreamStackBusLane[25][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane13_strm1_ready         ( DownstreamStackBusLane[25][13].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane13_strm1_cntl          ( DownstreamStackBusLane[25][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane13_strm1_data          ( DownstreamStackBusLane[25][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane13_strm1_data_valid    ( DownstreamStackBusLane[25][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane14_strm0_ready         ( DownstreamStackBusLane[25][14].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane14_strm0_cntl          ( DownstreamStackBusLane[25][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane14_strm0_data          ( DownstreamStackBusLane[25][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane14_strm0_data_valid    ( DownstreamStackBusLane[25][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane14_strm1_ready         ( DownstreamStackBusLane[25][14].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane14_strm1_cntl          ( DownstreamStackBusLane[25][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane14_strm1_data          ( DownstreamStackBusLane[25][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane14_strm1_data_valid    ( DownstreamStackBusLane[25][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane15_strm0_ready         ( DownstreamStackBusLane[25][15].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane15_strm0_cntl          ( DownstreamStackBusLane[25][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane15_strm0_data          ( DownstreamStackBusLane[25][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane15_strm0_data_valid    ( DownstreamStackBusLane[25][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane15_strm1_ready         ( DownstreamStackBusLane[25][15].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane15_strm1_cntl          ( DownstreamStackBusLane[25][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane15_strm1_data          ( DownstreamStackBusLane[25][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane15_strm1_data_valid    ( DownstreamStackBusLane[25][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane16_strm0_ready         ( DownstreamStackBusLane[25][16].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane16_strm0_cntl          ( DownstreamStackBusLane[25][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane16_strm0_data          ( DownstreamStackBusLane[25][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane16_strm0_data_valid    ( DownstreamStackBusLane[25][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane16_strm1_ready         ( DownstreamStackBusLane[25][16].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane16_strm1_cntl          ( DownstreamStackBusLane[25][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane16_strm1_data          ( DownstreamStackBusLane[25][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane16_strm1_data_valid    ( DownstreamStackBusLane[25][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane17_strm0_ready         ( DownstreamStackBusLane[25][17].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane17_strm0_cntl          ( DownstreamStackBusLane[25][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane17_strm0_data          ( DownstreamStackBusLane[25][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane17_strm0_data_valid    ( DownstreamStackBusLane[25][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane17_strm1_ready         ( DownstreamStackBusLane[25][17].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane17_strm1_cntl          ( DownstreamStackBusLane[25][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane17_strm1_data          ( DownstreamStackBusLane[25][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane17_strm1_data_valid    ( DownstreamStackBusLane[25][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane18_strm0_ready         ( DownstreamStackBusLane[25][18].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane18_strm0_cntl          ( DownstreamStackBusLane[25][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane18_strm0_data          ( DownstreamStackBusLane[25][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane18_strm0_data_valid    ( DownstreamStackBusLane[25][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane18_strm1_ready         ( DownstreamStackBusLane[25][18].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane18_strm1_cntl          ( DownstreamStackBusLane[25][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane18_strm1_data          ( DownstreamStackBusLane[25][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane18_strm1_data_valid    ( DownstreamStackBusLane[25][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane19_strm0_ready         ( DownstreamStackBusLane[25][19].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane19_strm0_cntl          ( DownstreamStackBusLane[25][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane19_strm0_data          ( DownstreamStackBusLane[25][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane19_strm0_data_valid    ( DownstreamStackBusLane[25][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane19_strm1_ready         ( DownstreamStackBusLane[25][19].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane19_strm1_cntl          ( DownstreamStackBusLane[25][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane19_strm1_data          ( DownstreamStackBusLane[25][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane19_strm1_data_valid    ( DownstreamStackBusLane[25][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane20_strm0_ready         ( DownstreamStackBusLane[25][20].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane20_strm0_cntl          ( DownstreamStackBusLane[25][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane20_strm0_data          ( DownstreamStackBusLane[25][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane20_strm0_data_valid    ( DownstreamStackBusLane[25][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane20_strm1_ready         ( DownstreamStackBusLane[25][20].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane20_strm1_cntl          ( DownstreamStackBusLane[25][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane20_strm1_data          ( DownstreamStackBusLane[25][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane20_strm1_data_valid    ( DownstreamStackBusLane[25][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane21_strm0_ready         ( DownstreamStackBusLane[25][21].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane21_strm0_cntl          ( DownstreamStackBusLane[25][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane21_strm0_data          ( DownstreamStackBusLane[25][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane21_strm0_data_valid    ( DownstreamStackBusLane[25][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane21_strm1_ready         ( DownstreamStackBusLane[25][21].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane21_strm1_cntl          ( DownstreamStackBusLane[25][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane21_strm1_data          ( DownstreamStackBusLane[25][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane21_strm1_data_valid    ( DownstreamStackBusLane[25][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane22_strm0_ready         ( DownstreamStackBusLane[25][22].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane22_strm0_cntl          ( DownstreamStackBusLane[25][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane22_strm0_data          ( DownstreamStackBusLane[25][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane22_strm0_data_valid    ( DownstreamStackBusLane[25][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane22_strm1_ready         ( DownstreamStackBusLane[25][22].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane22_strm1_cntl          ( DownstreamStackBusLane[25][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane22_strm1_data          ( DownstreamStackBusLane[25][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane22_strm1_data_valid    ( DownstreamStackBusLane[25][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane23_strm0_ready         ( DownstreamStackBusLane[25][23].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane23_strm0_cntl          ( DownstreamStackBusLane[25][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane23_strm0_data          ( DownstreamStackBusLane[25][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane23_strm0_data_valid    ( DownstreamStackBusLane[25][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane23_strm1_ready         ( DownstreamStackBusLane[25][23].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane23_strm1_cntl          ( DownstreamStackBusLane[25][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane23_strm1_data          ( DownstreamStackBusLane[25][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane23_strm1_data_valid    ( DownstreamStackBusLane[25][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane24_strm0_ready         ( DownstreamStackBusLane[25][24].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane24_strm0_cntl          ( DownstreamStackBusLane[25][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane24_strm0_data          ( DownstreamStackBusLane[25][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane24_strm0_data_valid    ( DownstreamStackBusLane[25][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane24_strm1_ready         ( DownstreamStackBusLane[25][24].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane24_strm1_cntl          ( DownstreamStackBusLane[25][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane24_strm1_data          ( DownstreamStackBusLane[25][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane24_strm1_data_valid    ( DownstreamStackBusLane[25][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane25_strm0_ready         ( DownstreamStackBusLane[25][25].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane25_strm0_cntl          ( DownstreamStackBusLane[25][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane25_strm0_data          ( DownstreamStackBusLane[25][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane25_strm0_data_valid    ( DownstreamStackBusLane[25][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane25_strm1_ready         ( DownstreamStackBusLane[25][25].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane25_strm1_cntl          ( DownstreamStackBusLane[25][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane25_strm1_data          ( DownstreamStackBusLane[25][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane25_strm1_data_valid    ( DownstreamStackBusLane[25][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane26_strm0_ready         ( DownstreamStackBusLane[25][26].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane26_strm0_cntl          ( DownstreamStackBusLane[25][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane26_strm0_data          ( DownstreamStackBusLane[25][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane26_strm0_data_valid    ( DownstreamStackBusLane[25][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane26_strm1_ready         ( DownstreamStackBusLane[25][26].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane26_strm1_cntl          ( DownstreamStackBusLane[25][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane26_strm1_data          ( DownstreamStackBusLane[25][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane26_strm1_data_valid    ( DownstreamStackBusLane[25][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane27_strm0_ready         ( DownstreamStackBusLane[25][27].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane27_strm0_cntl          ( DownstreamStackBusLane[25][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane27_strm0_data          ( DownstreamStackBusLane[25][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane27_strm0_data_valid    ( DownstreamStackBusLane[25][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane27_strm1_ready         ( DownstreamStackBusLane[25][27].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane27_strm1_cntl          ( DownstreamStackBusLane[25][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane27_strm1_data          ( DownstreamStackBusLane[25][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane27_strm1_data_valid    ( DownstreamStackBusLane[25][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane28_strm0_ready         ( DownstreamStackBusLane[25][28].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane28_strm0_cntl          ( DownstreamStackBusLane[25][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane28_strm0_data          ( DownstreamStackBusLane[25][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane28_strm0_data_valid    ( DownstreamStackBusLane[25][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane28_strm1_ready         ( DownstreamStackBusLane[25][28].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane28_strm1_cntl          ( DownstreamStackBusLane[25][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane28_strm1_data          ( DownstreamStackBusLane[25][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane28_strm1_data_valid    ( DownstreamStackBusLane[25][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane29_strm0_ready         ( DownstreamStackBusLane[25][29].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane29_strm0_cntl          ( DownstreamStackBusLane[25][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane29_strm0_data          ( DownstreamStackBusLane[25][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane29_strm0_data_valid    ( DownstreamStackBusLane[25][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane29_strm1_ready         ( DownstreamStackBusLane[25][29].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane29_strm1_cntl          ( DownstreamStackBusLane[25][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane29_strm1_data          ( DownstreamStackBusLane[25][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane29_strm1_data_valid    ( DownstreamStackBusLane[25][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane30_strm0_ready         ( DownstreamStackBusLane[25][30].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane30_strm0_cntl          ( DownstreamStackBusLane[25][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane30_strm0_data          ( DownstreamStackBusLane[25][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane30_strm0_data_valid    ( DownstreamStackBusLane[25][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane30_strm1_ready         ( DownstreamStackBusLane[25][30].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane30_strm1_cntl          ( DownstreamStackBusLane[25][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane30_strm1_data          ( DownstreamStackBusLane[25][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane30_strm1_data_valid    ( DownstreamStackBusLane[25][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 25, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane31_strm0_ready         ( DownstreamStackBusLane[25][31].pe__std__lane_strm0_ready              ),      
        .std__pe25__lane31_strm0_cntl          ( DownstreamStackBusLane[25][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe25__lane31_strm0_data          ( DownstreamStackBusLane[25][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe25__lane31_strm0_data_valid    ( DownstreamStackBusLane[25][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__std__lane31_strm1_ready         ( DownstreamStackBusLane[25][31].pe__std__lane_strm1_ready              ),      
        .std__pe25__lane31_strm1_cntl          ( DownstreamStackBusLane[25][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe25__lane31_strm1_data          ( DownstreamStackBusLane[25][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe25__lane31_strm1_data_valid    ( DownstreamStackBusLane[25][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane0_strm0_ready         ( DownstreamStackBusLane[26][0].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane0_strm0_cntl          ( DownstreamStackBusLane[26][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane0_strm0_data          ( DownstreamStackBusLane[26][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane0_strm0_data_valid    ( DownstreamStackBusLane[26][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane0_strm1_ready         ( DownstreamStackBusLane[26][0].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane0_strm1_cntl          ( DownstreamStackBusLane[26][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane0_strm1_data          ( DownstreamStackBusLane[26][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane0_strm1_data_valid    ( DownstreamStackBusLane[26][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane1_strm0_ready         ( DownstreamStackBusLane[26][1].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane1_strm0_cntl          ( DownstreamStackBusLane[26][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane1_strm0_data          ( DownstreamStackBusLane[26][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane1_strm0_data_valid    ( DownstreamStackBusLane[26][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane1_strm1_ready         ( DownstreamStackBusLane[26][1].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane1_strm1_cntl          ( DownstreamStackBusLane[26][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane1_strm1_data          ( DownstreamStackBusLane[26][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane1_strm1_data_valid    ( DownstreamStackBusLane[26][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane2_strm0_ready         ( DownstreamStackBusLane[26][2].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane2_strm0_cntl          ( DownstreamStackBusLane[26][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane2_strm0_data          ( DownstreamStackBusLane[26][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane2_strm0_data_valid    ( DownstreamStackBusLane[26][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane2_strm1_ready         ( DownstreamStackBusLane[26][2].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane2_strm1_cntl          ( DownstreamStackBusLane[26][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane2_strm1_data          ( DownstreamStackBusLane[26][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane2_strm1_data_valid    ( DownstreamStackBusLane[26][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane3_strm0_ready         ( DownstreamStackBusLane[26][3].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane3_strm0_cntl          ( DownstreamStackBusLane[26][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane3_strm0_data          ( DownstreamStackBusLane[26][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane3_strm0_data_valid    ( DownstreamStackBusLane[26][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane3_strm1_ready         ( DownstreamStackBusLane[26][3].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane3_strm1_cntl          ( DownstreamStackBusLane[26][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane3_strm1_data          ( DownstreamStackBusLane[26][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane3_strm1_data_valid    ( DownstreamStackBusLane[26][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane4_strm0_ready         ( DownstreamStackBusLane[26][4].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane4_strm0_cntl          ( DownstreamStackBusLane[26][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane4_strm0_data          ( DownstreamStackBusLane[26][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane4_strm0_data_valid    ( DownstreamStackBusLane[26][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane4_strm1_ready         ( DownstreamStackBusLane[26][4].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane4_strm1_cntl          ( DownstreamStackBusLane[26][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane4_strm1_data          ( DownstreamStackBusLane[26][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane4_strm1_data_valid    ( DownstreamStackBusLane[26][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane5_strm0_ready         ( DownstreamStackBusLane[26][5].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane5_strm0_cntl          ( DownstreamStackBusLane[26][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane5_strm0_data          ( DownstreamStackBusLane[26][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane5_strm0_data_valid    ( DownstreamStackBusLane[26][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane5_strm1_ready         ( DownstreamStackBusLane[26][5].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane5_strm1_cntl          ( DownstreamStackBusLane[26][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane5_strm1_data          ( DownstreamStackBusLane[26][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane5_strm1_data_valid    ( DownstreamStackBusLane[26][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane6_strm0_ready         ( DownstreamStackBusLane[26][6].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane6_strm0_cntl          ( DownstreamStackBusLane[26][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane6_strm0_data          ( DownstreamStackBusLane[26][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane6_strm0_data_valid    ( DownstreamStackBusLane[26][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane6_strm1_ready         ( DownstreamStackBusLane[26][6].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane6_strm1_cntl          ( DownstreamStackBusLane[26][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane6_strm1_data          ( DownstreamStackBusLane[26][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane6_strm1_data_valid    ( DownstreamStackBusLane[26][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane7_strm0_ready         ( DownstreamStackBusLane[26][7].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane7_strm0_cntl          ( DownstreamStackBusLane[26][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane7_strm0_data          ( DownstreamStackBusLane[26][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane7_strm0_data_valid    ( DownstreamStackBusLane[26][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane7_strm1_ready         ( DownstreamStackBusLane[26][7].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane7_strm1_cntl          ( DownstreamStackBusLane[26][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane7_strm1_data          ( DownstreamStackBusLane[26][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane7_strm1_data_valid    ( DownstreamStackBusLane[26][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane8_strm0_ready         ( DownstreamStackBusLane[26][8].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane8_strm0_cntl          ( DownstreamStackBusLane[26][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane8_strm0_data          ( DownstreamStackBusLane[26][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane8_strm0_data_valid    ( DownstreamStackBusLane[26][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane8_strm1_ready         ( DownstreamStackBusLane[26][8].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane8_strm1_cntl          ( DownstreamStackBusLane[26][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane8_strm1_data          ( DownstreamStackBusLane[26][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane8_strm1_data_valid    ( DownstreamStackBusLane[26][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane9_strm0_ready         ( DownstreamStackBusLane[26][9].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane9_strm0_cntl          ( DownstreamStackBusLane[26][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane9_strm0_data          ( DownstreamStackBusLane[26][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane9_strm0_data_valid    ( DownstreamStackBusLane[26][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane9_strm1_ready         ( DownstreamStackBusLane[26][9].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane9_strm1_cntl          ( DownstreamStackBusLane[26][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane9_strm1_data          ( DownstreamStackBusLane[26][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane9_strm1_data_valid    ( DownstreamStackBusLane[26][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane10_strm0_ready         ( DownstreamStackBusLane[26][10].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane10_strm0_cntl          ( DownstreamStackBusLane[26][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane10_strm0_data          ( DownstreamStackBusLane[26][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane10_strm0_data_valid    ( DownstreamStackBusLane[26][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane10_strm1_ready         ( DownstreamStackBusLane[26][10].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane10_strm1_cntl          ( DownstreamStackBusLane[26][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane10_strm1_data          ( DownstreamStackBusLane[26][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane10_strm1_data_valid    ( DownstreamStackBusLane[26][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane11_strm0_ready         ( DownstreamStackBusLane[26][11].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane11_strm0_cntl          ( DownstreamStackBusLane[26][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane11_strm0_data          ( DownstreamStackBusLane[26][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane11_strm0_data_valid    ( DownstreamStackBusLane[26][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane11_strm1_ready         ( DownstreamStackBusLane[26][11].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane11_strm1_cntl          ( DownstreamStackBusLane[26][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane11_strm1_data          ( DownstreamStackBusLane[26][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane11_strm1_data_valid    ( DownstreamStackBusLane[26][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane12_strm0_ready         ( DownstreamStackBusLane[26][12].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane12_strm0_cntl          ( DownstreamStackBusLane[26][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane12_strm0_data          ( DownstreamStackBusLane[26][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane12_strm0_data_valid    ( DownstreamStackBusLane[26][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane12_strm1_ready         ( DownstreamStackBusLane[26][12].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane12_strm1_cntl          ( DownstreamStackBusLane[26][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane12_strm1_data          ( DownstreamStackBusLane[26][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane12_strm1_data_valid    ( DownstreamStackBusLane[26][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane13_strm0_ready         ( DownstreamStackBusLane[26][13].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane13_strm0_cntl          ( DownstreamStackBusLane[26][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane13_strm0_data          ( DownstreamStackBusLane[26][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane13_strm0_data_valid    ( DownstreamStackBusLane[26][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane13_strm1_ready         ( DownstreamStackBusLane[26][13].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane13_strm1_cntl          ( DownstreamStackBusLane[26][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane13_strm1_data          ( DownstreamStackBusLane[26][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane13_strm1_data_valid    ( DownstreamStackBusLane[26][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane14_strm0_ready         ( DownstreamStackBusLane[26][14].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane14_strm0_cntl          ( DownstreamStackBusLane[26][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane14_strm0_data          ( DownstreamStackBusLane[26][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane14_strm0_data_valid    ( DownstreamStackBusLane[26][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane14_strm1_ready         ( DownstreamStackBusLane[26][14].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane14_strm1_cntl          ( DownstreamStackBusLane[26][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane14_strm1_data          ( DownstreamStackBusLane[26][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane14_strm1_data_valid    ( DownstreamStackBusLane[26][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane15_strm0_ready         ( DownstreamStackBusLane[26][15].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane15_strm0_cntl          ( DownstreamStackBusLane[26][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane15_strm0_data          ( DownstreamStackBusLane[26][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane15_strm0_data_valid    ( DownstreamStackBusLane[26][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane15_strm1_ready         ( DownstreamStackBusLane[26][15].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane15_strm1_cntl          ( DownstreamStackBusLane[26][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane15_strm1_data          ( DownstreamStackBusLane[26][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane15_strm1_data_valid    ( DownstreamStackBusLane[26][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane16_strm0_ready         ( DownstreamStackBusLane[26][16].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane16_strm0_cntl          ( DownstreamStackBusLane[26][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane16_strm0_data          ( DownstreamStackBusLane[26][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane16_strm0_data_valid    ( DownstreamStackBusLane[26][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane16_strm1_ready         ( DownstreamStackBusLane[26][16].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane16_strm1_cntl          ( DownstreamStackBusLane[26][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane16_strm1_data          ( DownstreamStackBusLane[26][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane16_strm1_data_valid    ( DownstreamStackBusLane[26][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane17_strm0_ready         ( DownstreamStackBusLane[26][17].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane17_strm0_cntl          ( DownstreamStackBusLane[26][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane17_strm0_data          ( DownstreamStackBusLane[26][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane17_strm0_data_valid    ( DownstreamStackBusLane[26][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane17_strm1_ready         ( DownstreamStackBusLane[26][17].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane17_strm1_cntl          ( DownstreamStackBusLane[26][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane17_strm1_data          ( DownstreamStackBusLane[26][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane17_strm1_data_valid    ( DownstreamStackBusLane[26][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane18_strm0_ready         ( DownstreamStackBusLane[26][18].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane18_strm0_cntl          ( DownstreamStackBusLane[26][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane18_strm0_data          ( DownstreamStackBusLane[26][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane18_strm0_data_valid    ( DownstreamStackBusLane[26][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane18_strm1_ready         ( DownstreamStackBusLane[26][18].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane18_strm1_cntl          ( DownstreamStackBusLane[26][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane18_strm1_data          ( DownstreamStackBusLane[26][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane18_strm1_data_valid    ( DownstreamStackBusLane[26][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane19_strm0_ready         ( DownstreamStackBusLane[26][19].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane19_strm0_cntl          ( DownstreamStackBusLane[26][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane19_strm0_data          ( DownstreamStackBusLane[26][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane19_strm0_data_valid    ( DownstreamStackBusLane[26][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane19_strm1_ready         ( DownstreamStackBusLane[26][19].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane19_strm1_cntl          ( DownstreamStackBusLane[26][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane19_strm1_data          ( DownstreamStackBusLane[26][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane19_strm1_data_valid    ( DownstreamStackBusLane[26][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane20_strm0_ready         ( DownstreamStackBusLane[26][20].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane20_strm0_cntl          ( DownstreamStackBusLane[26][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane20_strm0_data          ( DownstreamStackBusLane[26][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane20_strm0_data_valid    ( DownstreamStackBusLane[26][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane20_strm1_ready         ( DownstreamStackBusLane[26][20].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane20_strm1_cntl          ( DownstreamStackBusLane[26][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane20_strm1_data          ( DownstreamStackBusLane[26][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane20_strm1_data_valid    ( DownstreamStackBusLane[26][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane21_strm0_ready         ( DownstreamStackBusLane[26][21].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane21_strm0_cntl          ( DownstreamStackBusLane[26][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane21_strm0_data          ( DownstreamStackBusLane[26][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane21_strm0_data_valid    ( DownstreamStackBusLane[26][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane21_strm1_ready         ( DownstreamStackBusLane[26][21].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane21_strm1_cntl          ( DownstreamStackBusLane[26][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane21_strm1_data          ( DownstreamStackBusLane[26][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane21_strm1_data_valid    ( DownstreamStackBusLane[26][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane22_strm0_ready         ( DownstreamStackBusLane[26][22].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane22_strm0_cntl          ( DownstreamStackBusLane[26][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane22_strm0_data          ( DownstreamStackBusLane[26][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane22_strm0_data_valid    ( DownstreamStackBusLane[26][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane22_strm1_ready         ( DownstreamStackBusLane[26][22].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane22_strm1_cntl          ( DownstreamStackBusLane[26][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane22_strm1_data          ( DownstreamStackBusLane[26][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane22_strm1_data_valid    ( DownstreamStackBusLane[26][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane23_strm0_ready         ( DownstreamStackBusLane[26][23].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane23_strm0_cntl          ( DownstreamStackBusLane[26][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane23_strm0_data          ( DownstreamStackBusLane[26][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane23_strm0_data_valid    ( DownstreamStackBusLane[26][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane23_strm1_ready         ( DownstreamStackBusLane[26][23].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane23_strm1_cntl          ( DownstreamStackBusLane[26][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane23_strm1_data          ( DownstreamStackBusLane[26][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane23_strm1_data_valid    ( DownstreamStackBusLane[26][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane24_strm0_ready         ( DownstreamStackBusLane[26][24].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane24_strm0_cntl          ( DownstreamStackBusLane[26][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane24_strm0_data          ( DownstreamStackBusLane[26][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane24_strm0_data_valid    ( DownstreamStackBusLane[26][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane24_strm1_ready         ( DownstreamStackBusLane[26][24].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane24_strm1_cntl          ( DownstreamStackBusLane[26][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane24_strm1_data          ( DownstreamStackBusLane[26][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane24_strm1_data_valid    ( DownstreamStackBusLane[26][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane25_strm0_ready         ( DownstreamStackBusLane[26][25].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane25_strm0_cntl          ( DownstreamStackBusLane[26][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane25_strm0_data          ( DownstreamStackBusLane[26][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane25_strm0_data_valid    ( DownstreamStackBusLane[26][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane25_strm1_ready         ( DownstreamStackBusLane[26][25].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane25_strm1_cntl          ( DownstreamStackBusLane[26][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane25_strm1_data          ( DownstreamStackBusLane[26][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane25_strm1_data_valid    ( DownstreamStackBusLane[26][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane26_strm0_ready         ( DownstreamStackBusLane[26][26].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane26_strm0_cntl          ( DownstreamStackBusLane[26][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane26_strm0_data          ( DownstreamStackBusLane[26][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane26_strm0_data_valid    ( DownstreamStackBusLane[26][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane26_strm1_ready         ( DownstreamStackBusLane[26][26].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane26_strm1_cntl          ( DownstreamStackBusLane[26][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane26_strm1_data          ( DownstreamStackBusLane[26][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane26_strm1_data_valid    ( DownstreamStackBusLane[26][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane27_strm0_ready         ( DownstreamStackBusLane[26][27].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane27_strm0_cntl          ( DownstreamStackBusLane[26][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane27_strm0_data          ( DownstreamStackBusLane[26][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane27_strm0_data_valid    ( DownstreamStackBusLane[26][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane27_strm1_ready         ( DownstreamStackBusLane[26][27].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane27_strm1_cntl          ( DownstreamStackBusLane[26][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane27_strm1_data          ( DownstreamStackBusLane[26][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane27_strm1_data_valid    ( DownstreamStackBusLane[26][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane28_strm0_ready         ( DownstreamStackBusLane[26][28].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane28_strm0_cntl          ( DownstreamStackBusLane[26][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane28_strm0_data          ( DownstreamStackBusLane[26][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane28_strm0_data_valid    ( DownstreamStackBusLane[26][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane28_strm1_ready         ( DownstreamStackBusLane[26][28].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane28_strm1_cntl          ( DownstreamStackBusLane[26][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane28_strm1_data          ( DownstreamStackBusLane[26][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane28_strm1_data_valid    ( DownstreamStackBusLane[26][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane29_strm0_ready         ( DownstreamStackBusLane[26][29].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane29_strm0_cntl          ( DownstreamStackBusLane[26][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane29_strm0_data          ( DownstreamStackBusLane[26][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane29_strm0_data_valid    ( DownstreamStackBusLane[26][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane29_strm1_ready         ( DownstreamStackBusLane[26][29].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane29_strm1_cntl          ( DownstreamStackBusLane[26][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane29_strm1_data          ( DownstreamStackBusLane[26][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane29_strm1_data_valid    ( DownstreamStackBusLane[26][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane30_strm0_ready         ( DownstreamStackBusLane[26][30].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane30_strm0_cntl          ( DownstreamStackBusLane[26][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane30_strm0_data          ( DownstreamStackBusLane[26][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane30_strm0_data_valid    ( DownstreamStackBusLane[26][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane30_strm1_ready         ( DownstreamStackBusLane[26][30].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane30_strm1_cntl          ( DownstreamStackBusLane[26][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane30_strm1_data          ( DownstreamStackBusLane[26][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane30_strm1_data_valid    ( DownstreamStackBusLane[26][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 26, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane31_strm0_ready         ( DownstreamStackBusLane[26][31].pe__std__lane_strm0_ready              ),      
        .std__pe26__lane31_strm0_cntl          ( DownstreamStackBusLane[26][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe26__lane31_strm0_data          ( DownstreamStackBusLane[26][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe26__lane31_strm0_data_valid    ( DownstreamStackBusLane[26][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__std__lane31_strm1_ready         ( DownstreamStackBusLane[26][31].pe__std__lane_strm1_ready              ),      
        .std__pe26__lane31_strm1_cntl          ( DownstreamStackBusLane[26][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe26__lane31_strm1_data          ( DownstreamStackBusLane[26][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe26__lane31_strm1_data_valid    ( DownstreamStackBusLane[26][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane0_strm0_ready         ( DownstreamStackBusLane[27][0].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane0_strm0_cntl          ( DownstreamStackBusLane[27][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane0_strm0_data          ( DownstreamStackBusLane[27][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane0_strm0_data_valid    ( DownstreamStackBusLane[27][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane0_strm1_ready         ( DownstreamStackBusLane[27][0].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane0_strm1_cntl          ( DownstreamStackBusLane[27][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane0_strm1_data          ( DownstreamStackBusLane[27][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane0_strm1_data_valid    ( DownstreamStackBusLane[27][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane1_strm0_ready         ( DownstreamStackBusLane[27][1].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane1_strm0_cntl          ( DownstreamStackBusLane[27][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane1_strm0_data          ( DownstreamStackBusLane[27][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane1_strm0_data_valid    ( DownstreamStackBusLane[27][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane1_strm1_ready         ( DownstreamStackBusLane[27][1].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane1_strm1_cntl          ( DownstreamStackBusLane[27][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane1_strm1_data          ( DownstreamStackBusLane[27][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane1_strm1_data_valid    ( DownstreamStackBusLane[27][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane2_strm0_ready         ( DownstreamStackBusLane[27][2].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane2_strm0_cntl          ( DownstreamStackBusLane[27][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane2_strm0_data          ( DownstreamStackBusLane[27][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane2_strm0_data_valid    ( DownstreamStackBusLane[27][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane2_strm1_ready         ( DownstreamStackBusLane[27][2].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane2_strm1_cntl          ( DownstreamStackBusLane[27][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane2_strm1_data          ( DownstreamStackBusLane[27][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane2_strm1_data_valid    ( DownstreamStackBusLane[27][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane3_strm0_ready         ( DownstreamStackBusLane[27][3].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane3_strm0_cntl          ( DownstreamStackBusLane[27][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane3_strm0_data          ( DownstreamStackBusLane[27][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane3_strm0_data_valid    ( DownstreamStackBusLane[27][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane3_strm1_ready         ( DownstreamStackBusLane[27][3].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane3_strm1_cntl          ( DownstreamStackBusLane[27][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane3_strm1_data          ( DownstreamStackBusLane[27][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane3_strm1_data_valid    ( DownstreamStackBusLane[27][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane4_strm0_ready         ( DownstreamStackBusLane[27][4].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane4_strm0_cntl          ( DownstreamStackBusLane[27][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane4_strm0_data          ( DownstreamStackBusLane[27][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane4_strm0_data_valid    ( DownstreamStackBusLane[27][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane4_strm1_ready         ( DownstreamStackBusLane[27][4].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane4_strm1_cntl          ( DownstreamStackBusLane[27][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane4_strm1_data          ( DownstreamStackBusLane[27][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane4_strm1_data_valid    ( DownstreamStackBusLane[27][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane5_strm0_ready         ( DownstreamStackBusLane[27][5].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane5_strm0_cntl          ( DownstreamStackBusLane[27][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane5_strm0_data          ( DownstreamStackBusLane[27][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane5_strm0_data_valid    ( DownstreamStackBusLane[27][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane5_strm1_ready         ( DownstreamStackBusLane[27][5].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane5_strm1_cntl          ( DownstreamStackBusLane[27][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane5_strm1_data          ( DownstreamStackBusLane[27][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane5_strm1_data_valid    ( DownstreamStackBusLane[27][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane6_strm0_ready         ( DownstreamStackBusLane[27][6].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane6_strm0_cntl          ( DownstreamStackBusLane[27][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane6_strm0_data          ( DownstreamStackBusLane[27][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane6_strm0_data_valid    ( DownstreamStackBusLane[27][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane6_strm1_ready         ( DownstreamStackBusLane[27][6].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane6_strm1_cntl          ( DownstreamStackBusLane[27][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane6_strm1_data          ( DownstreamStackBusLane[27][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane6_strm1_data_valid    ( DownstreamStackBusLane[27][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane7_strm0_ready         ( DownstreamStackBusLane[27][7].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane7_strm0_cntl          ( DownstreamStackBusLane[27][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane7_strm0_data          ( DownstreamStackBusLane[27][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane7_strm0_data_valid    ( DownstreamStackBusLane[27][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane7_strm1_ready         ( DownstreamStackBusLane[27][7].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane7_strm1_cntl          ( DownstreamStackBusLane[27][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane7_strm1_data          ( DownstreamStackBusLane[27][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane7_strm1_data_valid    ( DownstreamStackBusLane[27][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane8_strm0_ready         ( DownstreamStackBusLane[27][8].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane8_strm0_cntl          ( DownstreamStackBusLane[27][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane8_strm0_data          ( DownstreamStackBusLane[27][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane8_strm0_data_valid    ( DownstreamStackBusLane[27][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane8_strm1_ready         ( DownstreamStackBusLane[27][8].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane8_strm1_cntl          ( DownstreamStackBusLane[27][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane8_strm1_data          ( DownstreamStackBusLane[27][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane8_strm1_data_valid    ( DownstreamStackBusLane[27][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane9_strm0_ready         ( DownstreamStackBusLane[27][9].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane9_strm0_cntl          ( DownstreamStackBusLane[27][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane9_strm0_data          ( DownstreamStackBusLane[27][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane9_strm0_data_valid    ( DownstreamStackBusLane[27][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane9_strm1_ready         ( DownstreamStackBusLane[27][9].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane9_strm1_cntl          ( DownstreamStackBusLane[27][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane9_strm1_data          ( DownstreamStackBusLane[27][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane9_strm1_data_valid    ( DownstreamStackBusLane[27][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane10_strm0_ready         ( DownstreamStackBusLane[27][10].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane10_strm0_cntl          ( DownstreamStackBusLane[27][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane10_strm0_data          ( DownstreamStackBusLane[27][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane10_strm0_data_valid    ( DownstreamStackBusLane[27][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane10_strm1_ready         ( DownstreamStackBusLane[27][10].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane10_strm1_cntl          ( DownstreamStackBusLane[27][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane10_strm1_data          ( DownstreamStackBusLane[27][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane10_strm1_data_valid    ( DownstreamStackBusLane[27][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane11_strm0_ready         ( DownstreamStackBusLane[27][11].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane11_strm0_cntl          ( DownstreamStackBusLane[27][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane11_strm0_data          ( DownstreamStackBusLane[27][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane11_strm0_data_valid    ( DownstreamStackBusLane[27][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane11_strm1_ready         ( DownstreamStackBusLane[27][11].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane11_strm1_cntl          ( DownstreamStackBusLane[27][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane11_strm1_data          ( DownstreamStackBusLane[27][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane11_strm1_data_valid    ( DownstreamStackBusLane[27][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane12_strm0_ready         ( DownstreamStackBusLane[27][12].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane12_strm0_cntl          ( DownstreamStackBusLane[27][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane12_strm0_data          ( DownstreamStackBusLane[27][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane12_strm0_data_valid    ( DownstreamStackBusLane[27][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane12_strm1_ready         ( DownstreamStackBusLane[27][12].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane12_strm1_cntl          ( DownstreamStackBusLane[27][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane12_strm1_data          ( DownstreamStackBusLane[27][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane12_strm1_data_valid    ( DownstreamStackBusLane[27][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane13_strm0_ready         ( DownstreamStackBusLane[27][13].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane13_strm0_cntl          ( DownstreamStackBusLane[27][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane13_strm0_data          ( DownstreamStackBusLane[27][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane13_strm0_data_valid    ( DownstreamStackBusLane[27][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane13_strm1_ready         ( DownstreamStackBusLane[27][13].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane13_strm1_cntl          ( DownstreamStackBusLane[27][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane13_strm1_data          ( DownstreamStackBusLane[27][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane13_strm1_data_valid    ( DownstreamStackBusLane[27][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane14_strm0_ready         ( DownstreamStackBusLane[27][14].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane14_strm0_cntl          ( DownstreamStackBusLane[27][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane14_strm0_data          ( DownstreamStackBusLane[27][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane14_strm0_data_valid    ( DownstreamStackBusLane[27][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane14_strm1_ready         ( DownstreamStackBusLane[27][14].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane14_strm1_cntl          ( DownstreamStackBusLane[27][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane14_strm1_data          ( DownstreamStackBusLane[27][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane14_strm1_data_valid    ( DownstreamStackBusLane[27][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane15_strm0_ready         ( DownstreamStackBusLane[27][15].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane15_strm0_cntl          ( DownstreamStackBusLane[27][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane15_strm0_data          ( DownstreamStackBusLane[27][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane15_strm0_data_valid    ( DownstreamStackBusLane[27][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane15_strm1_ready         ( DownstreamStackBusLane[27][15].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane15_strm1_cntl          ( DownstreamStackBusLane[27][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane15_strm1_data          ( DownstreamStackBusLane[27][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane15_strm1_data_valid    ( DownstreamStackBusLane[27][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane16_strm0_ready         ( DownstreamStackBusLane[27][16].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane16_strm0_cntl          ( DownstreamStackBusLane[27][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane16_strm0_data          ( DownstreamStackBusLane[27][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane16_strm0_data_valid    ( DownstreamStackBusLane[27][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane16_strm1_ready         ( DownstreamStackBusLane[27][16].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane16_strm1_cntl          ( DownstreamStackBusLane[27][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane16_strm1_data          ( DownstreamStackBusLane[27][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane16_strm1_data_valid    ( DownstreamStackBusLane[27][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane17_strm0_ready         ( DownstreamStackBusLane[27][17].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane17_strm0_cntl          ( DownstreamStackBusLane[27][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane17_strm0_data          ( DownstreamStackBusLane[27][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane17_strm0_data_valid    ( DownstreamStackBusLane[27][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane17_strm1_ready         ( DownstreamStackBusLane[27][17].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane17_strm1_cntl          ( DownstreamStackBusLane[27][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane17_strm1_data          ( DownstreamStackBusLane[27][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane17_strm1_data_valid    ( DownstreamStackBusLane[27][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane18_strm0_ready         ( DownstreamStackBusLane[27][18].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane18_strm0_cntl          ( DownstreamStackBusLane[27][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane18_strm0_data          ( DownstreamStackBusLane[27][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane18_strm0_data_valid    ( DownstreamStackBusLane[27][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane18_strm1_ready         ( DownstreamStackBusLane[27][18].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane18_strm1_cntl          ( DownstreamStackBusLane[27][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane18_strm1_data          ( DownstreamStackBusLane[27][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane18_strm1_data_valid    ( DownstreamStackBusLane[27][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane19_strm0_ready         ( DownstreamStackBusLane[27][19].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane19_strm0_cntl          ( DownstreamStackBusLane[27][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane19_strm0_data          ( DownstreamStackBusLane[27][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane19_strm0_data_valid    ( DownstreamStackBusLane[27][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane19_strm1_ready         ( DownstreamStackBusLane[27][19].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane19_strm1_cntl          ( DownstreamStackBusLane[27][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane19_strm1_data          ( DownstreamStackBusLane[27][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane19_strm1_data_valid    ( DownstreamStackBusLane[27][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane20_strm0_ready         ( DownstreamStackBusLane[27][20].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane20_strm0_cntl          ( DownstreamStackBusLane[27][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane20_strm0_data          ( DownstreamStackBusLane[27][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane20_strm0_data_valid    ( DownstreamStackBusLane[27][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane20_strm1_ready         ( DownstreamStackBusLane[27][20].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane20_strm1_cntl          ( DownstreamStackBusLane[27][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane20_strm1_data          ( DownstreamStackBusLane[27][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane20_strm1_data_valid    ( DownstreamStackBusLane[27][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane21_strm0_ready         ( DownstreamStackBusLane[27][21].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane21_strm0_cntl          ( DownstreamStackBusLane[27][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane21_strm0_data          ( DownstreamStackBusLane[27][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane21_strm0_data_valid    ( DownstreamStackBusLane[27][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane21_strm1_ready         ( DownstreamStackBusLane[27][21].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane21_strm1_cntl          ( DownstreamStackBusLane[27][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane21_strm1_data          ( DownstreamStackBusLane[27][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane21_strm1_data_valid    ( DownstreamStackBusLane[27][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane22_strm0_ready         ( DownstreamStackBusLane[27][22].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane22_strm0_cntl          ( DownstreamStackBusLane[27][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane22_strm0_data          ( DownstreamStackBusLane[27][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane22_strm0_data_valid    ( DownstreamStackBusLane[27][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane22_strm1_ready         ( DownstreamStackBusLane[27][22].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane22_strm1_cntl          ( DownstreamStackBusLane[27][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane22_strm1_data          ( DownstreamStackBusLane[27][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane22_strm1_data_valid    ( DownstreamStackBusLane[27][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane23_strm0_ready         ( DownstreamStackBusLane[27][23].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane23_strm0_cntl          ( DownstreamStackBusLane[27][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane23_strm0_data          ( DownstreamStackBusLane[27][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane23_strm0_data_valid    ( DownstreamStackBusLane[27][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane23_strm1_ready         ( DownstreamStackBusLane[27][23].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane23_strm1_cntl          ( DownstreamStackBusLane[27][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane23_strm1_data          ( DownstreamStackBusLane[27][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane23_strm1_data_valid    ( DownstreamStackBusLane[27][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane24_strm0_ready         ( DownstreamStackBusLane[27][24].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane24_strm0_cntl          ( DownstreamStackBusLane[27][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane24_strm0_data          ( DownstreamStackBusLane[27][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane24_strm0_data_valid    ( DownstreamStackBusLane[27][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane24_strm1_ready         ( DownstreamStackBusLane[27][24].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane24_strm1_cntl          ( DownstreamStackBusLane[27][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane24_strm1_data          ( DownstreamStackBusLane[27][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane24_strm1_data_valid    ( DownstreamStackBusLane[27][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane25_strm0_ready         ( DownstreamStackBusLane[27][25].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane25_strm0_cntl          ( DownstreamStackBusLane[27][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane25_strm0_data          ( DownstreamStackBusLane[27][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane25_strm0_data_valid    ( DownstreamStackBusLane[27][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane25_strm1_ready         ( DownstreamStackBusLane[27][25].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane25_strm1_cntl          ( DownstreamStackBusLane[27][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane25_strm1_data          ( DownstreamStackBusLane[27][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane25_strm1_data_valid    ( DownstreamStackBusLane[27][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane26_strm0_ready         ( DownstreamStackBusLane[27][26].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane26_strm0_cntl          ( DownstreamStackBusLane[27][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane26_strm0_data          ( DownstreamStackBusLane[27][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane26_strm0_data_valid    ( DownstreamStackBusLane[27][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane26_strm1_ready         ( DownstreamStackBusLane[27][26].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane26_strm1_cntl          ( DownstreamStackBusLane[27][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane26_strm1_data          ( DownstreamStackBusLane[27][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane26_strm1_data_valid    ( DownstreamStackBusLane[27][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane27_strm0_ready         ( DownstreamStackBusLane[27][27].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane27_strm0_cntl          ( DownstreamStackBusLane[27][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane27_strm0_data          ( DownstreamStackBusLane[27][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane27_strm0_data_valid    ( DownstreamStackBusLane[27][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane27_strm1_ready         ( DownstreamStackBusLane[27][27].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane27_strm1_cntl          ( DownstreamStackBusLane[27][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane27_strm1_data          ( DownstreamStackBusLane[27][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane27_strm1_data_valid    ( DownstreamStackBusLane[27][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane28_strm0_ready         ( DownstreamStackBusLane[27][28].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane28_strm0_cntl          ( DownstreamStackBusLane[27][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane28_strm0_data          ( DownstreamStackBusLane[27][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane28_strm0_data_valid    ( DownstreamStackBusLane[27][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane28_strm1_ready         ( DownstreamStackBusLane[27][28].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane28_strm1_cntl          ( DownstreamStackBusLane[27][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane28_strm1_data          ( DownstreamStackBusLane[27][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane28_strm1_data_valid    ( DownstreamStackBusLane[27][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane29_strm0_ready         ( DownstreamStackBusLane[27][29].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane29_strm0_cntl          ( DownstreamStackBusLane[27][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane29_strm0_data          ( DownstreamStackBusLane[27][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane29_strm0_data_valid    ( DownstreamStackBusLane[27][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane29_strm1_ready         ( DownstreamStackBusLane[27][29].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane29_strm1_cntl          ( DownstreamStackBusLane[27][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane29_strm1_data          ( DownstreamStackBusLane[27][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane29_strm1_data_valid    ( DownstreamStackBusLane[27][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane30_strm0_ready         ( DownstreamStackBusLane[27][30].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane30_strm0_cntl          ( DownstreamStackBusLane[27][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane30_strm0_data          ( DownstreamStackBusLane[27][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane30_strm0_data_valid    ( DownstreamStackBusLane[27][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane30_strm1_ready         ( DownstreamStackBusLane[27][30].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane30_strm1_cntl          ( DownstreamStackBusLane[27][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane30_strm1_data          ( DownstreamStackBusLane[27][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane30_strm1_data_valid    ( DownstreamStackBusLane[27][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 27, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane31_strm0_ready         ( DownstreamStackBusLane[27][31].pe__std__lane_strm0_ready              ),      
        .std__pe27__lane31_strm0_cntl          ( DownstreamStackBusLane[27][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe27__lane31_strm0_data          ( DownstreamStackBusLane[27][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe27__lane31_strm0_data_valid    ( DownstreamStackBusLane[27][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__std__lane31_strm1_ready         ( DownstreamStackBusLane[27][31].pe__std__lane_strm1_ready              ),      
        .std__pe27__lane31_strm1_cntl          ( DownstreamStackBusLane[27][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe27__lane31_strm1_data          ( DownstreamStackBusLane[27][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe27__lane31_strm1_data_valid    ( DownstreamStackBusLane[27][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane0_strm0_ready         ( DownstreamStackBusLane[28][0].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane0_strm0_cntl          ( DownstreamStackBusLane[28][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane0_strm0_data          ( DownstreamStackBusLane[28][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane0_strm0_data_valid    ( DownstreamStackBusLane[28][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane0_strm1_ready         ( DownstreamStackBusLane[28][0].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane0_strm1_cntl          ( DownstreamStackBusLane[28][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane0_strm1_data          ( DownstreamStackBusLane[28][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane0_strm1_data_valid    ( DownstreamStackBusLane[28][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane1_strm0_ready         ( DownstreamStackBusLane[28][1].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane1_strm0_cntl          ( DownstreamStackBusLane[28][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane1_strm0_data          ( DownstreamStackBusLane[28][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane1_strm0_data_valid    ( DownstreamStackBusLane[28][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane1_strm1_ready         ( DownstreamStackBusLane[28][1].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane1_strm1_cntl          ( DownstreamStackBusLane[28][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane1_strm1_data          ( DownstreamStackBusLane[28][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane1_strm1_data_valid    ( DownstreamStackBusLane[28][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane2_strm0_ready         ( DownstreamStackBusLane[28][2].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane2_strm0_cntl          ( DownstreamStackBusLane[28][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane2_strm0_data          ( DownstreamStackBusLane[28][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane2_strm0_data_valid    ( DownstreamStackBusLane[28][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane2_strm1_ready         ( DownstreamStackBusLane[28][2].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane2_strm1_cntl          ( DownstreamStackBusLane[28][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane2_strm1_data          ( DownstreamStackBusLane[28][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane2_strm1_data_valid    ( DownstreamStackBusLane[28][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane3_strm0_ready         ( DownstreamStackBusLane[28][3].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane3_strm0_cntl          ( DownstreamStackBusLane[28][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane3_strm0_data          ( DownstreamStackBusLane[28][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane3_strm0_data_valid    ( DownstreamStackBusLane[28][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane3_strm1_ready         ( DownstreamStackBusLane[28][3].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane3_strm1_cntl          ( DownstreamStackBusLane[28][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane3_strm1_data          ( DownstreamStackBusLane[28][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane3_strm1_data_valid    ( DownstreamStackBusLane[28][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane4_strm0_ready         ( DownstreamStackBusLane[28][4].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane4_strm0_cntl          ( DownstreamStackBusLane[28][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane4_strm0_data          ( DownstreamStackBusLane[28][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane4_strm0_data_valid    ( DownstreamStackBusLane[28][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane4_strm1_ready         ( DownstreamStackBusLane[28][4].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane4_strm1_cntl          ( DownstreamStackBusLane[28][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane4_strm1_data          ( DownstreamStackBusLane[28][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane4_strm1_data_valid    ( DownstreamStackBusLane[28][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane5_strm0_ready         ( DownstreamStackBusLane[28][5].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane5_strm0_cntl          ( DownstreamStackBusLane[28][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane5_strm0_data          ( DownstreamStackBusLane[28][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane5_strm0_data_valid    ( DownstreamStackBusLane[28][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane5_strm1_ready         ( DownstreamStackBusLane[28][5].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane5_strm1_cntl          ( DownstreamStackBusLane[28][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane5_strm1_data          ( DownstreamStackBusLane[28][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane5_strm1_data_valid    ( DownstreamStackBusLane[28][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane6_strm0_ready         ( DownstreamStackBusLane[28][6].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane6_strm0_cntl          ( DownstreamStackBusLane[28][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane6_strm0_data          ( DownstreamStackBusLane[28][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane6_strm0_data_valid    ( DownstreamStackBusLane[28][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane6_strm1_ready         ( DownstreamStackBusLane[28][6].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane6_strm1_cntl          ( DownstreamStackBusLane[28][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane6_strm1_data          ( DownstreamStackBusLane[28][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane6_strm1_data_valid    ( DownstreamStackBusLane[28][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane7_strm0_ready         ( DownstreamStackBusLane[28][7].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane7_strm0_cntl          ( DownstreamStackBusLane[28][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane7_strm0_data          ( DownstreamStackBusLane[28][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane7_strm0_data_valid    ( DownstreamStackBusLane[28][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane7_strm1_ready         ( DownstreamStackBusLane[28][7].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane7_strm1_cntl          ( DownstreamStackBusLane[28][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane7_strm1_data          ( DownstreamStackBusLane[28][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane7_strm1_data_valid    ( DownstreamStackBusLane[28][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane8_strm0_ready         ( DownstreamStackBusLane[28][8].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane8_strm0_cntl          ( DownstreamStackBusLane[28][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane8_strm0_data          ( DownstreamStackBusLane[28][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane8_strm0_data_valid    ( DownstreamStackBusLane[28][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane8_strm1_ready         ( DownstreamStackBusLane[28][8].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane8_strm1_cntl          ( DownstreamStackBusLane[28][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane8_strm1_data          ( DownstreamStackBusLane[28][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane8_strm1_data_valid    ( DownstreamStackBusLane[28][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane9_strm0_ready         ( DownstreamStackBusLane[28][9].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane9_strm0_cntl          ( DownstreamStackBusLane[28][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane9_strm0_data          ( DownstreamStackBusLane[28][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane9_strm0_data_valid    ( DownstreamStackBusLane[28][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane9_strm1_ready         ( DownstreamStackBusLane[28][9].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane9_strm1_cntl          ( DownstreamStackBusLane[28][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane9_strm1_data          ( DownstreamStackBusLane[28][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane9_strm1_data_valid    ( DownstreamStackBusLane[28][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane10_strm0_ready         ( DownstreamStackBusLane[28][10].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane10_strm0_cntl          ( DownstreamStackBusLane[28][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane10_strm0_data          ( DownstreamStackBusLane[28][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane10_strm0_data_valid    ( DownstreamStackBusLane[28][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane10_strm1_ready         ( DownstreamStackBusLane[28][10].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane10_strm1_cntl          ( DownstreamStackBusLane[28][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane10_strm1_data          ( DownstreamStackBusLane[28][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane10_strm1_data_valid    ( DownstreamStackBusLane[28][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane11_strm0_ready         ( DownstreamStackBusLane[28][11].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane11_strm0_cntl          ( DownstreamStackBusLane[28][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane11_strm0_data          ( DownstreamStackBusLane[28][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane11_strm0_data_valid    ( DownstreamStackBusLane[28][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane11_strm1_ready         ( DownstreamStackBusLane[28][11].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane11_strm1_cntl          ( DownstreamStackBusLane[28][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane11_strm1_data          ( DownstreamStackBusLane[28][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane11_strm1_data_valid    ( DownstreamStackBusLane[28][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane12_strm0_ready         ( DownstreamStackBusLane[28][12].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane12_strm0_cntl          ( DownstreamStackBusLane[28][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane12_strm0_data          ( DownstreamStackBusLane[28][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane12_strm0_data_valid    ( DownstreamStackBusLane[28][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane12_strm1_ready         ( DownstreamStackBusLane[28][12].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane12_strm1_cntl          ( DownstreamStackBusLane[28][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane12_strm1_data          ( DownstreamStackBusLane[28][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane12_strm1_data_valid    ( DownstreamStackBusLane[28][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane13_strm0_ready         ( DownstreamStackBusLane[28][13].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane13_strm0_cntl          ( DownstreamStackBusLane[28][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane13_strm0_data          ( DownstreamStackBusLane[28][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane13_strm0_data_valid    ( DownstreamStackBusLane[28][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane13_strm1_ready         ( DownstreamStackBusLane[28][13].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane13_strm1_cntl          ( DownstreamStackBusLane[28][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane13_strm1_data          ( DownstreamStackBusLane[28][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane13_strm1_data_valid    ( DownstreamStackBusLane[28][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane14_strm0_ready         ( DownstreamStackBusLane[28][14].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane14_strm0_cntl          ( DownstreamStackBusLane[28][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane14_strm0_data          ( DownstreamStackBusLane[28][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane14_strm0_data_valid    ( DownstreamStackBusLane[28][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane14_strm1_ready         ( DownstreamStackBusLane[28][14].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane14_strm1_cntl          ( DownstreamStackBusLane[28][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane14_strm1_data          ( DownstreamStackBusLane[28][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane14_strm1_data_valid    ( DownstreamStackBusLane[28][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane15_strm0_ready         ( DownstreamStackBusLane[28][15].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane15_strm0_cntl          ( DownstreamStackBusLane[28][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane15_strm0_data          ( DownstreamStackBusLane[28][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane15_strm0_data_valid    ( DownstreamStackBusLane[28][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane15_strm1_ready         ( DownstreamStackBusLane[28][15].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane15_strm1_cntl          ( DownstreamStackBusLane[28][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane15_strm1_data          ( DownstreamStackBusLane[28][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane15_strm1_data_valid    ( DownstreamStackBusLane[28][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane16_strm0_ready         ( DownstreamStackBusLane[28][16].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane16_strm0_cntl          ( DownstreamStackBusLane[28][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane16_strm0_data          ( DownstreamStackBusLane[28][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane16_strm0_data_valid    ( DownstreamStackBusLane[28][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane16_strm1_ready         ( DownstreamStackBusLane[28][16].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane16_strm1_cntl          ( DownstreamStackBusLane[28][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane16_strm1_data          ( DownstreamStackBusLane[28][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane16_strm1_data_valid    ( DownstreamStackBusLane[28][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane17_strm0_ready         ( DownstreamStackBusLane[28][17].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane17_strm0_cntl          ( DownstreamStackBusLane[28][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane17_strm0_data          ( DownstreamStackBusLane[28][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane17_strm0_data_valid    ( DownstreamStackBusLane[28][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane17_strm1_ready         ( DownstreamStackBusLane[28][17].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane17_strm1_cntl          ( DownstreamStackBusLane[28][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane17_strm1_data          ( DownstreamStackBusLane[28][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane17_strm1_data_valid    ( DownstreamStackBusLane[28][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane18_strm0_ready         ( DownstreamStackBusLane[28][18].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane18_strm0_cntl          ( DownstreamStackBusLane[28][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane18_strm0_data          ( DownstreamStackBusLane[28][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane18_strm0_data_valid    ( DownstreamStackBusLane[28][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane18_strm1_ready         ( DownstreamStackBusLane[28][18].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane18_strm1_cntl          ( DownstreamStackBusLane[28][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane18_strm1_data          ( DownstreamStackBusLane[28][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane18_strm1_data_valid    ( DownstreamStackBusLane[28][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane19_strm0_ready         ( DownstreamStackBusLane[28][19].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane19_strm0_cntl          ( DownstreamStackBusLane[28][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane19_strm0_data          ( DownstreamStackBusLane[28][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane19_strm0_data_valid    ( DownstreamStackBusLane[28][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane19_strm1_ready         ( DownstreamStackBusLane[28][19].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane19_strm1_cntl          ( DownstreamStackBusLane[28][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane19_strm1_data          ( DownstreamStackBusLane[28][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane19_strm1_data_valid    ( DownstreamStackBusLane[28][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane20_strm0_ready         ( DownstreamStackBusLane[28][20].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane20_strm0_cntl          ( DownstreamStackBusLane[28][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane20_strm0_data          ( DownstreamStackBusLane[28][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane20_strm0_data_valid    ( DownstreamStackBusLane[28][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane20_strm1_ready         ( DownstreamStackBusLane[28][20].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane20_strm1_cntl          ( DownstreamStackBusLane[28][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane20_strm1_data          ( DownstreamStackBusLane[28][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane20_strm1_data_valid    ( DownstreamStackBusLane[28][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane21_strm0_ready         ( DownstreamStackBusLane[28][21].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane21_strm0_cntl          ( DownstreamStackBusLane[28][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane21_strm0_data          ( DownstreamStackBusLane[28][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane21_strm0_data_valid    ( DownstreamStackBusLane[28][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane21_strm1_ready         ( DownstreamStackBusLane[28][21].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane21_strm1_cntl          ( DownstreamStackBusLane[28][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane21_strm1_data          ( DownstreamStackBusLane[28][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane21_strm1_data_valid    ( DownstreamStackBusLane[28][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane22_strm0_ready         ( DownstreamStackBusLane[28][22].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane22_strm0_cntl          ( DownstreamStackBusLane[28][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane22_strm0_data          ( DownstreamStackBusLane[28][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane22_strm0_data_valid    ( DownstreamStackBusLane[28][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane22_strm1_ready         ( DownstreamStackBusLane[28][22].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane22_strm1_cntl          ( DownstreamStackBusLane[28][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane22_strm1_data          ( DownstreamStackBusLane[28][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane22_strm1_data_valid    ( DownstreamStackBusLane[28][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane23_strm0_ready         ( DownstreamStackBusLane[28][23].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane23_strm0_cntl          ( DownstreamStackBusLane[28][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane23_strm0_data          ( DownstreamStackBusLane[28][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane23_strm0_data_valid    ( DownstreamStackBusLane[28][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane23_strm1_ready         ( DownstreamStackBusLane[28][23].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane23_strm1_cntl          ( DownstreamStackBusLane[28][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane23_strm1_data          ( DownstreamStackBusLane[28][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane23_strm1_data_valid    ( DownstreamStackBusLane[28][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane24_strm0_ready         ( DownstreamStackBusLane[28][24].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane24_strm0_cntl          ( DownstreamStackBusLane[28][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane24_strm0_data          ( DownstreamStackBusLane[28][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane24_strm0_data_valid    ( DownstreamStackBusLane[28][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane24_strm1_ready         ( DownstreamStackBusLane[28][24].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane24_strm1_cntl          ( DownstreamStackBusLane[28][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane24_strm1_data          ( DownstreamStackBusLane[28][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane24_strm1_data_valid    ( DownstreamStackBusLane[28][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane25_strm0_ready         ( DownstreamStackBusLane[28][25].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane25_strm0_cntl          ( DownstreamStackBusLane[28][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane25_strm0_data          ( DownstreamStackBusLane[28][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane25_strm0_data_valid    ( DownstreamStackBusLane[28][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane25_strm1_ready         ( DownstreamStackBusLane[28][25].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane25_strm1_cntl          ( DownstreamStackBusLane[28][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane25_strm1_data          ( DownstreamStackBusLane[28][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane25_strm1_data_valid    ( DownstreamStackBusLane[28][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane26_strm0_ready         ( DownstreamStackBusLane[28][26].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane26_strm0_cntl          ( DownstreamStackBusLane[28][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane26_strm0_data          ( DownstreamStackBusLane[28][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane26_strm0_data_valid    ( DownstreamStackBusLane[28][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane26_strm1_ready         ( DownstreamStackBusLane[28][26].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane26_strm1_cntl          ( DownstreamStackBusLane[28][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane26_strm1_data          ( DownstreamStackBusLane[28][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane26_strm1_data_valid    ( DownstreamStackBusLane[28][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane27_strm0_ready         ( DownstreamStackBusLane[28][27].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane27_strm0_cntl          ( DownstreamStackBusLane[28][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane27_strm0_data          ( DownstreamStackBusLane[28][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane27_strm0_data_valid    ( DownstreamStackBusLane[28][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane27_strm1_ready         ( DownstreamStackBusLane[28][27].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane27_strm1_cntl          ( DownstreamStackBusLane[28][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane27_strm1_data          ( DownstreamStackBusLane[28][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane27_strm1_data_valid    ( DownstreamStackBusLane[28][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane28_strm0_ready         ( DownstreamStackBusLane[28][28].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane28_strm0_cntl          ( DownstreamStackBusLane[28][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane28_strm0_data          ( DownstreamStackBusLane[28][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane28_strm0_data_valid    ( DownstreamStackBusLane[28][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane28_strm1_ready         ( DownstreamStackBusLane[28][28].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane28_strm1_cntl          ( DownstreamStackBusLane[28][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane28_strm1_data          ( DownstreamStackBusLane[28][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane28_strm1_data_valid    ( DownstreamStackBusLane[28][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane29_strm0_ready         ( DownstreamStackBusLane[28][29].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane29_strm0_cntl          ( DownstreamStackBusLane[28][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane29_strm0_data          ( DownstreamStackBusLane[28][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane29_strm0_data_valid    ( DownstreamStackBusLane[28][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane29_strm1_ready         ( DownstreamStackBusLane[28][29].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane29_strm1_cntl          ( DownstreamStackBusLane[28][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane29_strm1_data          ( DownstreamStackBusLane[28][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane29_strm1_data_valid    ( DownstreamStackBusLane[28][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane30_strm0_ready         ( DownstreamStackBusLane[28][30].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane30_strm0_cntl          ( DownstreamStackBusLane[28][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane30_strm0_data          ( DownstreamStackBusLane[28][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane30_strm0_data_valid    ( DownstreamStackBusLane[28][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane30_strm1_ready         ( DownstreamStackBusLane[28][30].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane30_strm1_cntl          ( DownstreamStackBusLane[28][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane30_strm1_data          ( DownstreamStackBusLane[28][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane30_strm1_data_valid    ( DownstreamStackBusLane[28][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 28, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane31_strm0_ready         ( DownstreamStackBusLane[28][31].pe__std__lane_strm0_ready              ),      
        .std__pe28__lane31_strm0_cntl          ( DownstreamStackBusLane[28][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe28__lane31_strm0_data          ( DownstreamStackBusLane[28][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe28__lane31_strm0_data_valid    ( DownstreamStackBusLane[28][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__std__lane31_strm1_ready         ( DownstreamStackBusLane[28][31].pe__std__lane_strm1_ready              ),      
        .std__pe28__lane31_strm1_cntl          ( DownstreamStackBusLane[28][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe28__lane31_strm1_data          ( DownstreamStackBusLane[28][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe28__lane31_strm1_data_valid    ( DownstreamStackBusLane[28][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane0_strm0_ready         ( DownstreamStackBusLane[29][0].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane0_strm0_cntl          ( DownstreamStackBusLane[29][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane0_strm0_data          ( DownstreamStackBusLane[29][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane0_strm0_data_valid    ( DownstreamStackBusLane[29][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane0_strm1_ready         ( DownstreamStackBusLane[29][0].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane0_strm1_cntl          ( DownstreamStackBusLane[29][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane0_strm1_data          ( DownstreamStackBusLane[29][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane0_strm1_data_valid    ( DownstreamStackBusLane[29][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane1_strm0_ready         ( DownstreamStackBusLane[29][1].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane1_strm0_cntl          ( DownstreamStackBusLane[29][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane1_strm0_data          ( DownstreamStackBusLane[29][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane1_strm0_data_valid    ( DownstreamStackBusLane[29][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane1_strm1_ready         ( DownstreamStackBusLane[29][1].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane1_strm1_cntl          ( DownstreamStackBusLane[29][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane1_strm1_data          ( DownstreamStackBusLane[29][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane1_strm1_data_valid    ( DownstreamStackBusLane[29][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane2_strm0_ready         ( DownstreamStackBusLane[29][2].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane2_strm0_cntl          ( DownstreamStackBusLane[29][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane2_strm0_data          ( DownstreamStackBusLane[29][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane2_strm0_data_valid    ( DownstreamStackBusLane[29][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane2_strm1_ready         ( DownstreamStackBusLane[29][2].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane2_strm1_cntl          ( DownstreamStackBusLane[29][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane2_strm1_data          ( DownstreamStackBusLane[29][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane2_strm1_data_valid    ( DownstreamStackBusLane[29][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane3_strm0_ready         ( DownstreamStackBusLane[29][3].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane3_strm0_cntl          ( DownstreamStackBusLane[29][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane3_strm0_data          ( DownstreamStackBusLane[29][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane3_strm0_data_valid    ( DownstreamStackBusLane[29][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane3_strm1_ready         ( DownstreamStackBusLane[29][3].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane3_strm1_cntl          ( DownstreamStackBusLane[29][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane3_strm1_data          ( DownstreamStackBusLane[29][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane3_strm1_data_valid    ( DownstreamStackBusLane[29][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane4_strm0_ready         ( DownstreamStackBusLane[29][4].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane4_strm0_cntl          ( DownstreamStackBusLane[29][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane4_strm0_data          ( DownstreamStackBusLane[29][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane4_strm0_data_valid    ( DownstreamStackBusLane[29][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane4_strm1_ready         ( DownstreamStackBusLane[29][4].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane4_strm1_cntl          ( DownstreamStackBusLane[29][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane4_strm1_data          ( DownstreamStackBusLane[29][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane4_strm1_data_valid    ( DownstreamStackBusLane[29][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane5_strm0_ready         ( DownstreamStackBusLane[29][5].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane5_strm0_cntl          ( DownstreamStackBusLane[29][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane5_strm0_data          ( DownstreamStackBusLane[29][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane5_strm0_data_valid    ( DownstreamStackBusLane[29][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane5_strm1_ready         ( DownstreamStackBusLane[29][5].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane5_strm1_cntl          ( DownstreamStackBusLane[29][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane5_strm1_data          ( DownstreamStackBusLane[29][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane5_strm1_data_valid    ( DownstreamStackBusLane[29][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane6_strm0_ready         ( DownstreamStackBusLane[29][6].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane6_strm0_cntl          ( DownstreamStackBusLane[29][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane6_strm0_data          ( DownstreamStackBusLane[29][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane6_strm0_data_valid    ( DownstreamStackBusLane[29][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane6_strm1_ready         ( DownstreamStackBusLane[29][6].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane6_strm1_cntl          ( DownstreamStackBusLane[29][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane6_strm1_data          ( DownstreamStackBusLane[29][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane6_strm1_data_valid    ( DownstreamStackBusLane[29][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane7_strm0_ready         ( DownstreamStackBusLane[29][7].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane7_strm0_cntl          ( DownstreamStackBusLane[29][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane7_strm0_data          ( DownstreamStackBusLane[29][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane7_strm0_data_valid    ( DownstreamStackBusLane[29][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane7_strm1_ready         ( DownstreamStackBusLane[29][7].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane7_strm1_cntl          ( DownstreamStackBusLane[29][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane7_strm1_data          ( DownstreamStackBusLane[29][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane7_strm1_data_valid    ( DownstreamStackBusLane[29][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane8_strm0_ready         ( DownstreamStackBusLane[29][8].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane8_strm0_cntl          ( DownstreamStackBusLane[29][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane8_strm0_data          ( DownstreamStackBusLane[29][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane8_strm0_data_valid    ( DownstreamStackBusLane[29][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane8_strm1_ready         ( DownstreamStackBusLane[29][8].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane8_strm1_cntl          ( DownstreamStackBusLane[29][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane8_strm1_data          ( DownstreamStackBusLane[29][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane8_strm1_data_valid    ( DownstreamStackBusLane[29][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane9_strm0_ready         ( DownstreamStackBusLane[29][9].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane9_strm0_cntl          ( DownstreamStackBusLane[29][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane9_strm0_data          ( DownstreamStackBusLane[29][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane9_strm0_data_valid    ( DownstreamStackBusLane[29][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane9_strm1_ready         ( DownstreamStackBusLane[29][9].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane9_strm1_cntl          ( DownstreamStackBusLane[29][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane9_strm1_data          ( DownstreamStackBusLane[29][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane9_strm1_data_valid    ( DownstreamStackBusLane[29][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane10_strm0_ready         ( DownstreamStackBusLane[29][10].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane10_strm0_cntl          ( DownstreamStackBusLane[29][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane10_strm0_data          ( DownstreamStackBusLane[29][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane10_strm0_data_valid    ( DownstreamStackBusLane[29][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane10_strm1_ready         ( DownstreamStackBusLane[29][10].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane10_strm1_cntl          ( DownstreamStackBusLane[29][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane10_strm1_data          ( DownstreamStackBusLane[29][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane10_strm1_data_valid    ( DownstreamStackBusLane[29][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane11_strm0_ready         ( DownstreamStackBusLane[29][11].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane11_strm0_cntl          ( DownstreamStackBusLane[29][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane11_strm0_data          ( DownstreamStackBusLane[29][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane11_strm0_data_valid    ( DownstreamStackBusLane[29][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane11_strm1_ready         ( DownstreamStackBusLane[29][11].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane11_strm1_cntl          ( DownstreamStackBusLane[29][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane11_strm1_data          ( DownstreamStackBusLane[29][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane11_strm1_data_valid    ( DownstreamStackBusLane[29][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane12_strm0_ready         ( DownstreamStackBusLane[29][12].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane12_strm0_cntl          ( DownstreamStackBusLane[29][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane12_strm0_data          ( DownstreamStackBusLane[29][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane12_strm0_data_valid    ( DownstreamStackBusLane[29][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane12_strm1_ready         ( DownstreamStackBusLane[29][12].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane12_strm1_cntl          ( DownstreamStackBusLane[29][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane12_strm1_data          ( DownstreamStackBusLane[29][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane12_strm1_data_valid    ( DownstreamStackBusLane[29][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane13_strm0_ready         ( DownstreamStackBusLane[29][13].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane13_strm0_cntl          ( DownstreamStackBusLane[29][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane13_strm0_data          ( DownstreamStackBusLane[29][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane13_strm0_data_valid    ( DownstreamStackBusLane[29][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane13_strm1_ready         ( DownstreamStackBusLane[29][13].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane13_strm1_cntl          ( DownstreamStackBusLane[29][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane13_strm1_data          ( DownstreamStackBusLane[29][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane13_strm1_data_valid    ( DownstreamStackBusLane[29][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane14_strm0_ready         ( DownstreamStackBusLane[29][14].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane14_strm0_cntl          ( DownstreamStackBusLane[29][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane14_strm0_data          ( DownstreamStackBusLane[29][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane14_strm0_data_valid    ( DownstreamStackBusLane[29][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane14_strm1_ready         ( DownstreamStackBusLane[29][14].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane14_strm1_cntl          ( DownstreamStackBusLane[29][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane14_strm1_data          ( DownstreamStackBusLane[29][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane14_strm1_data_valid    ( DownstreamStackBusLane[29][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane15_strm0_ready         ( DownstreamStackBusLane[29][15].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane15_strm0_cntl          ( DownstreamStackBusLane[29][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane15_strm0_data          ( DownstreamStackBusLane[29][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane15_strm0_data_valid    ( DownstreamStackBusLane[29][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane15_strm1_ready         ( DownstreamStackBusLane[29][15].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane15_strm1_cntl          ( DownstreamStackBusLane[29][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane15_strm1_data          ( DownstreamStackBusLane[29][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane15_strm1_data_valid    ( DownstreamStackBusLane[29][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane16_strm0_ready         ( DownstreamStackBusLane[29][16].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane16_strm0_cntl          ( DownstreamStackBusLane[29][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane16_strm0_data          ( DownstreamStackBusLane[29][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane16_strm0_data_valid    ( DownstreamStackBusLane[29][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane16_strm1_ready         ( DownstreamStackBusLane[29][16].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane16_strm1_cntl          ( DownstreamStackBusLane[29][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane16_strm1_data          ( DownstreamStackBusLane[29][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane16_strm1_data_valid    ( DownstreamStackBusLane[29][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane17_strm0_ready         ( DownstreamStackBusLane[29][17].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane17_strm0_cntl          ( DownstreamStackBusLane[29][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane17_strm0_data          ( DownstreamStackBusLane[29][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane17_strm0_data_valid    ( DownstreamStackBusLane[29][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane17_strm1_ready         ( DownstreamStackBusLane[29][17].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane17_strm1_cntl          ( DownstreamStackBusLane[29][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane17_strm1_data          ( DownstreamStackBusLane[29][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane17_strm1_data_valid    ( DownstreamStackBusLane[29][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane18_strm0_ready         ( DownstreamStackBusLane[29][18].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane18_strm0_cntl          ( DownstreamStackBusLane[29][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane18_strm0_data          ( DownstreamStackBusLane[29][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane18_strm0_data_valid    ( DownstreamStackBusLane[29][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane18_strm1_ready         ( DownstreamStackBusLane[29][18].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane18_strm1_cntl          ( DownstreamStackBusLane[29][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane18_strm1_data          ( DownstreamStackBusLane[29][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane18_strm1_data_valid    ( DownstreamStackBusLane[29][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane19_strm0_ready         ( DownstreamStackBusLane[29][19].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane19_strm0_cntl          ( DownstreamStackBusLane[29][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane19_strm0_data          ( DownstreamStackBusLane[29][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane19_strm0_data_valid    ( DownstreamStackBusLane[29][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane19_strm1_ready         ( DownstreamStackBusLane[29][19].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane19_strm1_cntl          ( DownstreamStackBusLane[29][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane19_strm1_data          ( DownstreamStackBusLane[29][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane19_strm1_data_valid    ( DownstreamStackBusLane[29][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane20_strm0_ready         ( DownstreamStackBusLane[29][20].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane20_strm0_cntl          ( DownstreamStackBusLane[29][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane20_strm0_data          ( DownstreamStackBusLane[29][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane20_strm0_data_valid    ( DownstreamStackBusLane[29][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane20_strm1_ready         ( DownstreamStackBusLane[29][20].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane20_strm1_cntl          ( DownstreamStackBusLane[29][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane20_strm1_data          ( DownstreamStackBusLane[29][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane20_strm1_data_valid    ( DownstreamStackBusLane[29][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane21_strm0_ready         ( DownstreamStackBusLane[29][21].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane21_strm0_cntl          ( DownstreamStackBusLane[29][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane21_strm0_data          ( DownstreamStackBusLane[29][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane21_strm0_data_valid    ( DownstreamStackBusLane[29][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane21_strm1_ready         ( DownstreamStackBusLane[29][21].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane21_strm1_cntl          ( DownstreamStackBusLane[29][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane21_strm1_data          ( DownstreamStackBusLane[29][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane21_strm1_data_valid    ( DownstreamStackBusLane[29][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane22_strm0_ready         ( DownstreamStackBusLane[29][22].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane22_strm0_cntl          ( DownstreamStackBusLane[29][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane22_strm0_data          ( DownstreamStackBusLane[29][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane22_strm0_data_valid    ( DownstreamStackBusLane[29][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane22_strm1_ready         ( DownstreamStackBusLane[29][22].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane22_strm1_cntl          ( DownstreamStackBusLane[29][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane22_strm1_data          ( DownstreamStackBusLane[29][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane22_strm1_data_valid    ( DownstreamStackBusLane[29][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane23_strm0_ready         ( DownstreamStackBusLane[29][23].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane23_strm0_cntl          ( DownstreamStackBusLane[29][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane23_strm0_data          ( DownstreamStackBusLane[29][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane23_strm0_data_valid    ( DownstreamStackBusLane[29][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane23_strm1_ready         ( DownstreamStackBusLane[29][23].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane23_strm1_cntl          ( DownstreamStackBusLane[29][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane23_strm1_data          ( DownstreamStackBusLane[29][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane23_strm1_data_valid    ( DownstreamStackBusLane[29][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane24_strm0_ready         ( DownstreamStackBusLane[29][24].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane24_strm0_cntl          ( DownstreamStackBusLane[29][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane24_strm0_data          ( DownstreamStackBusLane[29][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane24_strm0_data_valid    ( DownstreamStackBusLane[29][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane24_strm1_ready         ( DownstreamStackBusLane[29][24].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane24_strm1_cntl          ( DownstreamStackBusLane[29][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane24_strm1_data          ( DownstreamStackBusLane[29][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane24_strm1_data_valid    ( DownstreamStackBusLane[29][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane25_strm0_ready         ( DownstreamStackBusLane[29][25].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane25_strm0_cntl          ( DownstreamStackBusLane[29][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane25_strm0_data          ( DownstreamStackBusLane[29][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane25_strm0_data_valid    ( DownstreamStackBusLane[29][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane25_strm1_ready         ( DownstreamStackBusLane[29][25].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane25_strm1_cntl          ( DownstreamStackBusLane[29][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane25_strm1_data          ( DownstreamStackBusLane[29][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane25_strm1_data_valid    ( DownstreamStackBusLane[29][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane26_strm0_ready         ( DownstreamStackBusLane[29][26].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane26_strm0_cntl          ( DownstreamStackBusLane[29][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane26_strm0_data          ( DownstreamStackBusLane[29][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane26_strm0_data_valid    ( DownstreamStackBusLane[29][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane26_strm1_ready         ( DownstreamStackBusLane[29][26].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane26_strm1_cntl          ( DownstreamStackBusLane[29][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane26_strm1_data          ( DownstreamStackBusLane[29][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane26_strm1_data_valid    ( DownstreamStackBusLane[29][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane27_strm0_ready         ( DownstreamStackBusLane[29][27].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane27_strm0_cntl          ( DownstreamStackBusLane[29][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane27_strm0_data          ( DownstreamStackBusLane[29][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane27_strm0_data_valid    ( DownstreamStackBusLane[29][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane27_strm1_ready         ( DownstreamStackBusLane[29][27].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane27_strm1_cntl          ( DownstreamStackBusLane[29][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane27_strm1_data          ( DownstreamStackBusLane[29][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane27_strm1_data_valid    ( DownstreamStackBusLane[29][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane28_strm0_ready         ( DownstreamStackBusLane[29][28].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane28_strm0_cntl          ( DownstreamStackBusLane[29][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane28_strm0_data          ( DownstreamStackBusLane[29][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane28_strm0_data_valid    ( DownstreamStackBusLane[29][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane28_strm1_ready         ( DownstreamStackBusLane[29][28].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane28_strm1_cntl          ( DownstreamStackBusLane[29][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane28_strm1_data          ( DownstreamStackBusLane[29][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane28_strm1_data_valid    ( DownstreamStackBusLane[29][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane29_strm0_ready         ( DownstreamStackBusLane[29][29].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane29_strm0_cntl          ( DownstreamStackBusLane[29][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane29_strm0_data          ( DownstreamStackBusLane[29][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane29_strm0_data_valid    ( DownstreamStackBusLane[29][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane29_strm1_ready         ( DownstreamStackBusLane[29][29].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane29_strm1_cntl          ( DownstreamStackBusLane[29][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane29_strm1_data          ( DownstreamStackBusLane[29][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane29_strm1_data_valid    ( DownstreamStackBusLane[29][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane30_strm0_ready         ( DownstreamStackBusLane[29][30].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane30_strm0_cntl          ( DownstreamStackBusLane[29][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane30_strm0_data          ( DownstreamStackBusLane[29][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane30_strm0_data_valid    ( DownstreamStackBusLane[29][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane30_strm1_ready         ( DownstreamStackBusLane[29][30].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane30_strm1_cntl          ( DownstreamStackBusLane[29][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane30_strm1_data          ( DownstreamStackBusLane[29][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane30_strm1_data_valid    ( DownstreamStackBusLane[29][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 29, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane31_strm0_ready         ( DownstreamStackBusLane[29][31].pe__std__lane_strm0_ready              ),      
        .std__pe29__lane31_strm0_cntl          ( DownstreamStackBusLane[29][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe29__lane31_strm0_data          ( DownstreamStackBusLane[29][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe29__lane31_strm0_data_valid    ( DownstreamStackBusLane[29][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__std__lane31_strm1_ready         ( DownstreamStackBusLane[29][31].pe__std__lane_strm1_ready              ),      
        .std__pe29__lane31_strm1_cntl          ( DownstreamStackBusLane[29][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe29__lane31_strm1_data          ( DownstreamStackBusLane[29][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe29__lane31_strm1_data_valid    ( DownstreamStackBusLane[29][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane0_strm0_ready         ( DownstreamStackBusLane[30][0].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane0_strm0_cntl          ( DownstreamStackBusLane[30][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane0_strm0_data          ( DownstreamStackBusLane[30][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane0_strm0_data_valid    ( DownstreamStackBusLane[30][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane0_strm1_ready         ( DownstreamStackBusLane[30][0].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane0_strm1_cntl          ( DownstreamStackBusLane[30][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane0_strm1_data          ( DownstreamStackBusLane[30][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane0_strm1_data_valid    ( DownstreamStackBusLane[30][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane1_strm0_ready         ( DownstreamStackBusLane[30][1].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane1_strm0_cntl          ( DownstreamStackBusLane[30][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane1_strm0_data          ( DownstreamStackBusLane[30][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane1_strm0_data_valid    ( DownstreamStackBusLane[30][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane1_strm1_ready         ( DownstreamStackBusLane[30][1].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane1_strm1_cntl          ( DownstreamStackBusLane[30][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane1_strm1_data          ( DownstreamStackBusLane[30][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane1_strm1_data_valid    ( DownstreamStackBusLane[30][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane2_strm0_ready         ( DownstreamStackBusLane[30][2].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane2_strm0_cntl          ( DownstreamStackBusLane[30][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane2_strm0_data          ( DownstreamStackBusLane[30][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane2_strm0_data_valid    ( DownstreamStackBusLane[30][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane2_strm1_ready         ( DownstreamStackBusLane[30][2].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane2_strm1_cntl          ( DownstreamStackBusLane[30][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane2_strm1_data          ( DownstreamStackBusLane[30][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane2_strm1_data_valid    ( DownstreamStackBusLane[30][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane3_strm0_ready         ( DownstreamStackBusLane[30][3].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane3_strm0_cntl          ( DownstreamStackBusLane[30][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane3_strm0_data          ( DownstreamStackBusLane[30][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane3_strm0_data_valid    ( DownstreamStackBusLane[30][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane3_strm1_ready         ( DownstreamStackBusLane[30][3].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane3_strm1_cntl          ( DownstreamStackBusLane[30][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane3_strm1_data          ( DownstreamStackBusLane[30][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane3_strm1_data_valid    ( DownstreamStackBusLane[30][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane4_strm0_ready         ( DownstreamStackBusLane[30][4].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane4_strm0_cntl          ( DownstreamStackBusLane[30][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane4_strm0_data          ( DownstreamStackBusLane[30][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane4_strm0_data_valid    ( DownstreamStackBusLane[30][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane4_strm1_ready         ( DownstreamStackBusLane[30][4].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane4_strm1_cntl          ( DownstreamStackBusLane[30][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane4_strm1_data          ( DownstreamStackBusLane[30][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane4_strm1_data_valid    ( DownstreamStackBusLane[30][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane5_strm0_ready         ( DownstreamStackBusLane[30][5].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane5_strm0_cntl          ( DownstreamStackBusLane[30][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane5_strm0_data          ( DownstreamStackBusLane[30][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane5_strm0_data_valid    ( DownstreamStackBusLane[30][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane5_strm1_ready         ( DownstreamStackBusLane[30][5].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane5_strm1_cntl          ( DownstreamStackBusLane[30][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane5_strm1_data          ( DownstreamStackBusLane[30][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane5_strm1_data_valid    ( DownstreamStackBusLane[30][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane6_strm0_ready         ( DownstreamStackBusLane[30][6].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane6_strm0_cntl          ( DownstreamStackBusLane[30][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane6_strm0_data          ( DownstreamStackBusLane[30][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane6_strm0_data_valid    ( DownstreamStackBusLane[30][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane6_strm1_ready         ( DownstreamStackBusLane[30][6].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane6_strm1_cntl          ( DownstreamStackBusLane[30][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane6_strm1_data          ( DownstreamStackBusLane[30][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane6_strm1_data_valid    ( DownstreamStackBusLane[30][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane7_strm0_ready         ( DownstreamStackBusLane[30][7].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane7_strm0_cntl          ( DownstreamStackBusLane[30][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane7_strm0_data          ( DownstreamStackBusLane[30][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane7_strm0_data_valid    ( DownstreamStackBusLane[30][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane7_strm1_ready         ( DownstreamStackBusLane[30][7].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane7_strm1_cntl          ( DownstreamStackBusLane[30][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane7_strm1_data          ( DownstreamStackBusLane[30][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane7_strm1_data_valid    ( DownstreamStackBusLane[30][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane8_strm0_ready         ( DownstreamStackBusLane[30][8].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane8_strm0_cntl          ( DownstreamStackBusLane[30][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane8_strm0_data          ( DownstreamStackBusLane[30][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane8_strm0_data_valid    ( DownstreamStackBusLane[30][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane8_strm1_ready         ( DownstreamStackBusLane[30][8].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane8_strm1_cntl          ( DownstreamStackBusLane[30][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane8_strm1_data          ( DownstreamStackBusLane[30][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane8_strm1_data_valid    ( DownstreamStackBusLane[30][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane9_strm0_ready         ( DownstreamStackBusLane[30][9].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane9_strm0_cntl          ( DownstreamStackBusLane[30][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane9_strm0_data          ( DownstreamStackBusLane[30][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane9_strm0_data_valid    ( DownstreamStackBusLane[30][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane9_strm1_ready         ( DownstreamStackBusLane[30][9].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane9_strm1_cntl          ( DownstreamStackBusLane[30][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane9_strm1_data          ( DownstreamStackBusLane[30][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane9_strm1_data_valid    ( DownstreamStackBusLane[30][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane10_strm0_ready         ( DownstreamStackBusLane[30][10].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane10_strm0_cntl          ( DownstreamStackBusLane[30][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane10_strm0_data          ( DownstreamStackBusLane[30][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane10_strm0_data_valid    ( DownstreamStackBusLane[30][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane10_strm1_ready         ( DownstreamStackBusLane[30][10].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane10_strm1_cntl          ( DownstreamStackBusLane[30][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane10_strm1_data          ( DownstreamStackBusLane[30][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane10_strm1_data_valid    ( DownstreamStackBusLane[30][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane11_strm0_ready         ( DownstreamStackBusLane[30][11].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane11_strm0_cntl          ( DownstreamStackBusLane[30][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane11_strm0_data          ( DownstreamStackBusLane[30][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane11_strm0_data_valid    ( DownstreamStackBusLane[30][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane11_strm1_ready         ( DownstreamStackBusLane[30][11].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane11_strm1_cntl          ( DownstreamStackBusLane[30][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane11_strm1_data          ( DownstreamStackBusLane[30][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane11_strm1_data_valid    ( DownstreamStackBusLane[30][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane12_strm0_ready         ( DownstreamStackBusLane[30][12].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane12_strm0_cntl          ( DownstreamStackBusLane[30][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane12_strm0_data          ( DownstreamStackBusLane[30][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane12_strm0_data_valid    ( DownstreamStackBusLane[30][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane12_strm1_ready         ( DownstreamStackBusLane[30][12].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane12_strm1_cntl          ( DownstreamStackBusLane[30][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane12_strm1_data          ( DownstreamStackBusLane[30][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane12_strm1_data_valid    ( DownstreamStackBusLane[30][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane13_strm0_ready         ( DownstreamStackBusLane[30][13].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane13_strm0_cntl          ( DownstreamStackBusLane[30][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane13_strm0_data          ( DownstreamStackBusLane[30][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane13_strm0_data_valid    ( DownstreamStackBusLane[30][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane13_strm1_ready         ( DownstreamStackBusLane[30][13].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane13_strm1_cntl          ( DownstreamStackBusLane[30][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane13_strm1_data          ( DownstreamStackBusLane[30][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane13_strm1_data_valid    ( DownstreamStackBusLane[30][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane14_strm0_ready         ( DownstreamStackBusLane[30][14].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane14_strm0_cntl          ( DownstreamStackBusLane[30][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane14_strm0_data          ( DownstreamStackBusLane[30][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane14_strm0_data_valid    ( DownstreamStackBusLane[30][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane14_strm1_ready         ( DownstreamStackBusLane[30][14].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane14_strm1_cntl          ( DownstreamStackBusLane[30][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane14_strm1_data          ( DownstreamStackBusLane[30][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane14_strm1_data_valid    ( DownstreamStackBusLane[30][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane15_strm0_ready         ( DownstreamStackBusLane[30][15].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane15_strm0_cntl          ( DownstreamStackBusLane[30][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane15_strm0_data          ( DownstreamStackBusLane[30][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane15_strm0_data_valid    ( DownstreamStackBusLane[30][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane15_strm1_ready         ( DownstreamStackBusLane[30][15].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane15_strm1_cntl          ( DownstreamStackBusLane[30][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane15_strm1_data          ( DownstreamStackBusLane[30][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane15_strm1_data_valid    ( DownstreamStackBusLane[30][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane16_strm0_ready         ( DownstreamStackBusLane[30][16].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane16_strm0_cntl          ( DownstreamStackBusLane[30][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane16_strm0_data          ( DownstreamStackBusLane[30][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane16_strm0_data_valid    ( DownstreamStackBusLane[30][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane16_strm1_ready         ( DownstreamStackBusLane[30][16].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane16_strm1_cntl          ( DownstreamStackBusLane[30][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane16_strm1_data          ( DownstreamStackBusLane[30][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane16_strm1_data_valid    ( DownstreamStackBusLane[30][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane17_strm0_ready         ( DownstreamStackBusLane[30][17].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane17_strm0_cntl          ( DownstreamStackBusLane[30][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane17_strm0_data          ( DownstreamStackBusLane[30][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane17_strm0_data_valid    ( DownstreamStackBusLane[30][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane17_strm1_ready         ( DownstreamStackBusLane[30][17].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane17_strm1_cntl          ( DownstreamStackBusLane[30][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane17_strm1_data          ( DownstreamStackBusLane[30][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane17_strm1_data_valid    ( DownstreamStackBusLane[30][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane18_strm0_ready         ( DownstreamStackBusLane[30][18].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane18_strm0_cntl          ( DownstreamStackBusLane[30][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane18_strm0_data          ( DownstreamStackBusLane[30][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane18_strm0_data_valid    ( DownstreamStackBusLane[30][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane18_strm1_ready         ( DownstreamStackBusLane[30][18].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane18_strm1_cntl          ( DownstreamStackBusLane[30][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane18_strm1_data          ( DownstreamStackBusLane[30][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane18_strm1_data_valid    ( DownstreamStackBusLane[30][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane19_strm0_ready         ( DownstreamStackBusLane[30][19].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane19_strm0_cntl          ( DownstreamStackBusLane[30][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane19_strm0_data          ( DownstreamStackBusLane[30][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane19_strm0_data_valid    ( DownstreamStackBusLane[30][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane19_strm1_ready         ( DownstreamStackBusLane[30][19].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane19_strm1_cntl          ( DownstreamStackBusLane[30][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane19_strm1_data          ( DownstreamStackBusLane[30][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane19_strm1_data_valid    ( DownstreamStackBusLane[30][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane20_strm0_ready         ( DownstreamStackBusLane[30][20].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane20_strm0_cntl          ( DownstreamStackBusLane[30][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane20_strm0_data          ( DownstreamStackBusLane[30][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane20_strm0_data_valid    ( DownstreamStackBusLane[30][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane20_strm1_ready         ( DownstreamStackBusLane[30][20].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane20_strm1_cntl          ( DownstreamStackBusLane[30][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane20_strm1_data          ( DownstreamStackBusLane[30][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane20_strm1_data_valid    ( DownstreamStackBusLane[30][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane21_strm0_ready         ( DownstreamStackBusLane[30][21].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane21_strm0_cntl          ( DownstreamStackBusLane[30][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane21_strm0_data          ( DownstreamStackBusLane[30][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane21_strm0_data_valid    ( DownstreamStackBusLane[30][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane21_strm1_ready         ( DownstreamStackBusLane[30][21].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane21_strm1_cntl          ( DownstreamStackBusLane[30][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane21_strm1_data          ( DownstreamStackBusLane[30][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane21_strm1_data_valid    ( DownstreamStackBusLane[30][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane22_strm0_ready         ( DownstreamStackBusLane[30][22].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane22_strm0_cntl          ( DownstreamStackBusLane[30][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane22_strm0_data          ( DownstreamStackBusLane[30][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane22_strm0_data_valid    ( DownstreamStackBusLane[30][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane22_strm1_ready         ( DownstreamStackBusLane[30][22].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane22_strm1_cntl          ( DownstreamStackBusLane[30][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane22_strm1_data          ( DownstreamStackBusLane[30][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane22_strm1_data_valid    ( DownstreamStackBusLane[30][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane23_strm0_ready         ( DownstreamStackBusLane[30][23].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane23_strm0_cntl          ( DownstreamStackBusLane[30][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane23_strm0_data          ( DownstreamStackBusLane[30][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane23_strm0_data_valid    ( DownstreamStackBusLane[30][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane23_strm1_ready         ( DownstreamStackBusLane[30][23].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane23_strm1_cntl          ( DownstreamStackBusLane[30][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane23_strm1_data          ( DownstreamStackBusLane[30][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane23_strm1_data_valid    ( DownstreamStackBusLane[30][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane24_strm0_ready         ( DownstreamStackBusLane[30][24].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane24_strm0_cntl          ( DownstreamStackBusLane[30][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane24_strm0_data          ( DownstreamStackBusLane[30][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane24_strm0_data_valid    ( DownstreamStackBusLane[30][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane24_strm1_ready         ( DownstreamStackBusLane[30][24].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane24_strm1_cntl          ( DownstreamStackBusLane[30][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane24_strm1_data          ( DownstreamStackBusLane[30][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane24_strm1_data_valid    ( DownstreamStackBusLane[30][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane25_strm0_ready         ( DownstreamStackBusLane[30][25].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane25_strm0_cntl          ( DownstreamStackBusLane[30][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane25_strm0_data          ( DownstreamStackBusLane[30][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane25_strm0_data_valid    ( DownstreamStackBusLane[30][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane25_strm1_ready         ( DownstreamStackBusLane[30][25].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane25_strm1_cntl          ( DownstreamStackBusLane[30][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane25_strm1_data          ( DownstreamStackBusLane[30][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane25_strm1_data_valid    ( DownstreamStackBusLane[30][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane26_strm0_ready         ( DownstreamStackBusLane[30][26].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane26_strm0_cntl          ( DownstreamStackBusLane[30][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane26_strm0_data          ( DownstreamStackBusLane[30][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane26_strm0_data_valid    ( DownstreamStackBusLane[30][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane26_strm1_ready         ( DownstreamStackBusLane[30][26].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane26_strm1_cntl          ( DownstreamStackBusLane[30][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane26_strm1_data          ( DownstreamStackBusLane[30][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane26_strm1_data_valid    ( DownstreamStackBusLane[30][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane27_strm0_ready         ( DownstreamStackBusLane[30][27].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane27_strm0_cntl          ( DownstreamStackBusLane[30][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane27_strm0_data          ( DownstreamStackBusLane[30][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane27_strm0_data_valid    ( DownstreamStackBusLane[30][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane27_strm1_ready         ( DownstreamStackBusLane[30][27].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane27_strm1_cntl          ( DownstreamStackBusLane[30][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane27_strm1_data          ( DownstreamStackBusLane[30][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane27_strm1_data_valid    ( DownstreamStackBusLane[30][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane28_strm0_ready         ( DownstreamStackBusLane[30][28].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane28_strm0_cntl          ( DownstreamStackBusLane[30][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane28_strm0_data          ( DownstreamStackBusLane[30][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane28_strm0_data_valid    ( DownstreamStackBusLane[30][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane28_strm1_ready         ( DownstreamStackBusLane[30][28].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane28_strm1_cntl          ( DownstreamStackBusLane[30][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane28_strm1_data          ( DownstreamStackBusLane[30][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane28_strm1_data_valid    ( DownstreamStackBusLane[30][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane29_strm0_ready         ( DownstreamStackBusLane[30][29].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane29_strm0_cntl          ( DownstreamStackBusLane[30][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane29_strm0_data          ( DownstreamStackBusLane[30][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane29_strm0_data_valid    ( DownstreamStackBusLane[30][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane29_strm1_ready         ( DownstreamStackBusLane[30][29].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane29_strm1_cntl          ( DownstreamStackBusLane[30][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane29_strm1_data          ( DownstreamStackBusLane[30][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane29_strm1_data_valid    ( DownstreamStackBusLane[30][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane30_strm0_ready         ( DownstreamStackBusLane[30][30].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane30_strm0_cntl          ( DownstreamStackBusLane[30][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane30_strm0_data          ( DownstreamStackBusLane[30][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane30_strm0_data_valid    ( DownstreamStackBusLane[30][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane30_strm1_ready         ( DownstreamStackBusLane[30][30].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane30_strm1_cntl          ( DownstreamStackBusLane[30][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane30_strm1_data          ( DownstreamStackBusLane[30][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane30_strm1_data_valid    ( DownstreamStackBusLane[30][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 30, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane31_strm0_ready         ( DownstreamStackBusLane[30][31].pe__std__lane_strm0_ready              ),      
        .std__pe30__lane31_strm0_cntl          ( DownstreamStackBusLane[30][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe30__lane31_strm0_data          ( DownstreamStackBusLane[30][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe30__lane31_strm0_data_valid    ( DownstreamStackBusLane[30][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__std__lane31_strm1_ready         ( DownstreamStackBusLane[30][31].pe__std__lane_strm1_ready              ),      
        .std__pe30__lane31_strm1_cntl          ( DownstreamStackBusLane[30][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe30__lane31_strm1_data          ( DownstreamStackBusLane[30][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe30__lane31_strm1_data_valid    ( DownstreamStackBusLane[30][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane0_strm0_ready         ( DownstreamStackBusLane[31][0].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane0_strm0_cntl          ( DownstreamStackBusLane[31][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane0_strm0_data          ( DownstreamStackBusLane[31][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane0_strm0_data_valid    ( DownstreamStackBusLane[31][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane0_strm1_ready         ( DownstreamStackBusLane[31][0].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane0_strm1_cntl          ( DownstreamStackBusLane[31][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane0_strm1_data          ( DownstreamStackBusLane[31][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane0_strm1_data_valid    ( DownstreamStackBusLane[31][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane1_strm0_ready         ( DownstreamStackBusLane[31][1].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane1_strm0_cntl          ( DownstreamStackBusLane[31][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane1_strm0_data          ( DownstreamStackBusLane[31][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane1_strm0_data_valid    ( DownstreamStackBusLane[31][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane1_strm1_ready         ( DownstreamStackBusLane[31][1].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane1_strm1_cntl          ( DownstreamStackBusLane[31][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane1_strm1_data          ( DownstreamStackBusLane[31][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane1_strm1_data_valid    ( DownstreamStackBusLane[31][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane2_strm0_ready         ( DownstreamStackBusLane[31][2].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane2_strm0_cntl          ( DownstreamStackBusLane[31][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane2_strm0_data          ( DownstreamStackBusLane[31][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane2_strm0_data_valid    ( DownstreamStackBusLane[31][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane2_strm1_ready         ( DownstreamStackBusLane[31][2].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane2_strm1_cntl          ( DownstreamStackBusLane[31][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane2_strm1_data          ( DownstreamStackBusLane[31][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane2_strm1_data_valid    ( DownstreamStackBusLane[31][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane3_strm0_ready         ( DownstreamStackBusLane[31][3].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane3_strm0_cntl          ( DownstreamStackBusLane[31][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane3_strm0_data          ( DownstreamStackBusLane[31][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane3_strm0_data_valid    ( DownstreamStackBusLane[31][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane3_strm1_ready         ( DownstreamStackBusLane[31][3].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane3_strm1_cntl          ( DownstreamStackBusLane[31][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane3_strm1_data          ( DownstreamStackBusLane[31][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane3_strm1_data_valid    ( DownstreamStackBusLane[31][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane4_strm0_ready         ( DownstreamStackBusLane[31][4].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane4_strm0_cntl          ( DownstreamStackBusLane[31][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane4_strm0_data          ( DownstreamStackBusLane[31][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane4_strm0_data_valid    ( DownstreamStackBusLane[31][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane4_strm1_ready         ( DownstreamStackBusLane[31][4].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane4_strm1_cntl          ( DownstreamStackBusLane[31][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane4_strm1_data          ( DownstreamStackBusLane[31][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane4_strm1_data_valid    ( DownstreamStackBusLane[31][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane5_strm0_ready         ( DownstreamStackBusLane[31][5].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane5_strm0_cntl          ( DownstreamStackBusLane[31][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane5_strm0_data          ( DownstreamStackBusLane[31][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane5_strm0_data_valid    ( DownstreamStackBusLane[31][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane5_strm1_ready         ( DownstreamStackBusLane[31][5].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane5_strm1_cntl          ( DownstreamStackBusLane[31][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane5_strm1_data          ( DownstreamStackBusLane[31][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane5_strm1_data_valid    ( DownstreamStackBusLane[31][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane6_strm0_ready         ( DownstreamStackBusLane[31][6].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane6_strm0_cntl          ( DownstreamStackBusLane[31][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane6_strm0_data          ( DownstreamStackBusLane[31][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane6_strm0_data_valid    ( DownstreamStackBusLane[31][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane6_strm1_ready         ( DownstreamStackBusLane[31][6].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane6_strm1_cntl          ( DownstreamStackBusLane[31][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane6_strm1_data          ( DownstreamStackBusLane[31][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane6_strm1_data_valid    ( DownstreamStackBusLane[31][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane7_strm0_ready         ( DownstreamStackBusLane[31][7].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane7_strm0_cntl          ( DownstreamStackBusLane[31][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane7_strm0_data          ( DownstreamStackBusLane[31][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane7_strm0_data_valid    ( DownstreamStackBusLane[31][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane7_strm1_ready         ( DownstreamStackBusLane[31][7].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane7_strm1_cntl          ( DownstreamStackBusLane[31][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane7_strm1_data          ( DownstreamStackBusLane[31][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane7_strm1_data_valid    ( DownstreamStackBusLane[31][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane8_strm0_ready         ( DownstreamStackBusLane[31][8].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane8_strm0_cntl          ( DownstreamStackBusLane[31][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane8_strm0_data          ( DownstreamStackBusLane[31][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane8_strm0_data_valid    ( DownstreamStackBusLane[31][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane8_strm1_ready         ( DownstreamStackBusLane[31][8].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane8_strm1_cntl          ( DownstreamStackBusLane[31][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane8_strm1_data          ( DownstreamStackBusLane[31][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane8_strm1_data_valid    ( DownstreamStackBusLane[31][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane9_strm0_ready         ( DownstreamStackBusLane[31][9].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane9_strm0_cntl          ( DownstreamStackBusLane[31][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane9_strm0_data          ( DownstreamStackBusLane[31][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane9_strm0_data_valid    ( DownstreamStackBusLane[31][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane9_strm1_ready         ( DownstreamStackBusLane[31][9].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane9_strm1_cntl          ( DownstreamStackBusLane[31][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane9_strm1_data          ( DownstreamStackBusLane[31][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane9_strm1_data_valid    ( DownstreamStackBusLane[31][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane10_strm0_ready         ( DownstreamStackBusLane[31][10].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane10_strm0_cntl          ( DownstreamStackBusLane[31][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane10_strm0_data          ( DownstreamStackBusLane[31][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane10_strm0_data_valid    ( DownstreamStackBusLane[31][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane10_strm1_ready         ( DownstreamStackBusLane[31][10].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane10_strm1_cntl          ( DownstreamStackBusLane[31][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane10_strm1_data          ( DownstreamStackBusLane[31][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane10_strm1_data_valid    ( DownstreamStackBusLane[31][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane11_strm0_ready         ( DownstreamStackBusLane[31][11].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane11_strm0_cntl          ( DownstreamStackBusLane[31][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane11_strm0_data          ( DownstreamStackBusLane[31][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane11_strm0_data_valid    ( DownstreamStackBusLane[31][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane11_strm1_ready         ( DownstreamStackBusLane[31][11].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane11_strm1_cntl          ( DownstreamStackBusLane[31][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane11_strm1_data          ( DownstreamStackBusLane[31][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane11_strm1_data_valid    ( DownstreamStackBusLane[31][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane12_strm0_ready         ( DownstreamStackBusLane[31][12].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane12_strm0_cntl          ( DownstreamStackBusLane[31][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane12_strm0_data          ( DownstreamStackBusLane[31][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane12_strm0_data_valid    ( DownstreamStackBusLane[31][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane12_strm1_ready         ( DownstreamStackBusLane[31][12].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane12_strm1_cntl          ( DownstreamStackBusLane[31][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane12_strm1_data          ( DownstreamStackBusLane[31][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane12_strm1_data_valid    ( DownstreamStackBusLane[31][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane13_strm0_ready         ( DownstreamStackBusLane[31][13].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane13_strm0_cntl          ( DownstreamStackBusLane[31][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane13_strm0_data          ( DownstreamStackBusLane[31][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane13_strm0_data_valid    ( DownstreamStackBusLane[31][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane13_strm1_ready         ( DownstreamStackBusLane[31][13].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane13_strm1_cntl          ( DownstreamStackBusLane[31][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane13_strm1_data          ( DownstreamStackBusLane[31][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane13_strm1_data_valid    ( DownstreamStackBusLane[31][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane14_strm0_ready         ( DownstreamStackBusLane[31][14].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane14_strm0_cntl          ( DownstreamStackBusLane[31][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane14_strm0_data          ( DownstreamStackBusLane[31][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane14_strm0_data_valid    ( DownstreamStackBusLane[31][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane14_strm1_ready         ( DownstreamStackBusLane[31][14].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane14_strm1_cntl          ( DownstreamStackBusLane[31][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane14_strm1_data          ( DownstreamStackBusLane[31][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane14_strm1_data_valid    ( DownstreamStackBusLane[31][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane15_strm0_ready         ( DownstreamStackBusLane[31][15].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane15_strm0_cntl          ( DownstreamStackBusLane[31][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane15_strm0_data          ( DownstreamStackBusLane[31][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane15_strm0_data_valid    ( DownstreamStackBusLane[31][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane15_strm1_ready         ( DownstreamStackBusLane[31][15].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane15_strm1_cntl          ( DownstreamStackBusLane[31][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane15_strm1_data          ( DownstreamStackBusLane[31][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane15_strm1_data_valid    ( DownstreamStackBusLane[31][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane16_strm0_ready         ( DownstreamStackBusLane[31][16].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane16_strm0_cntl          ( DownstreamStackBusLane[31][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane16_strm0_data          ( DownstreamStackBusLane[31][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane16_strm0_data_valid    ( DownstreamStackBusLane[31][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane16_strm1_ready         ( DownstreamStackBusLane[31][16].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane16_strm1_cntl          ( DownstreamStackBusLane[31][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane16_strm1_data          ( DownstreamStackBusLane[31][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane16_strm1_data_valid    ( DownstreamStackBusLane[31][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane17_strm0_ready         ( DownstreamStackBusLane[31][17].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane17_strm0_cntl          ( DownstreamStackBusLane[31][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane17_strm0_data          ( DownstreamStackBusLane[31][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane17_strm0_data_valid    ( DownstreamStackBusLane[31][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane17_strm1_ready         ( DownstreamStackBusLane[31][17].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane17_strm1_cntl          ( DownstreamStackBusLane[31][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane17_strm1_data          ( DownstreamStackBusLane[31][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane17_strm1_data_valid    ( DownstreamStackBusLane[31][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane18_strm0_ready         ( DownstreamStackBusLane[31][18].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane18_strm0_cntl          ( DownstreamStackBusLane[31][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane18_strm0_data          ( DownstreamStackBusLane[31][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane18_strm0_data_valid    ( DownstreamStackBusLane[31][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane18_strm1_ready         ( DownstreamStackBusLane[31][18].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane18_strm1_cntl          ( DownstreamStackBusLane[31][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane18_strm1_data          ( DownstreamStackBusLane[31][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane18_strm1_data_valid    ( DownstreamStackBusLane[31][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane19_strm0_ready         ( DownstreamStackBusLane[31][19].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane19_strm0_cntl          ( DownstreamStackBusLane[31][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane19_strm0_data          ( DownstreamStackBusLane[31][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane19_strm0_data_valid    ( DownstreamStackBusLane[31][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane19_strm1_ready         ( DownstreamStackBusLane[31][19].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane19_strm1_cntl          ( DownstreamStackBusLane[31][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane19_strm1_data          ( DownstreamStackBusLane[31][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane19_strm1_data_valid    ( DownstreamStackBusLane[31][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane20_strm0_ready         ( DownstreamStackBusLane[31][20].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane20_strm0_cntl          ( DownstreamStackBusLane[31][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane20_strm0_data          ( DownstreamStackBusLane[31][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane20_strm0_data_valid    ( DownstreamStackBusLane[31][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane20_strm1_ready         ( DownstreamStackBusLane[31][20].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane20_strm1_cntl          ( DownstreamStackBusLane[31][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane20_strm1_data          ( DownstreamStackBusLane[31][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane20_strm1_data_valid    ( DownstreamStackBusLane[31][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane21_strm0_ready         ( DownstreamStackBusLane[31][21].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane21_strm0_cntl          ( DownstreamStackBusLane[31][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane21_strm0_data          ( DownstreamStackBusLane[31][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane21_strm0_data_valid    ( DownstreamStackBusLane[31][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane21_strm1_ready         ( DownstreamStackBusLane[31][21].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane21_strm1_cntl          ( DownstreamStackBusLane[31][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane21_strm1_data          ( DownstreamStackBusLane[31][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane21_strm1_data_valid    ( DownstreamStackBusLane[31][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane22_strm0_ready         ( DownstreamStackBusLane[31][22].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane22_strm0_cntl          ( DownstreamStackBusLane[31][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane22_strm0_data          ( DownstreamStackBusLane[31][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane22_strm0_data_valid    ( DownstreamStackBusLane[31][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane22_strm1_ready         ( DownstreamStackBusLane[31][22].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane22_strm1_cntl          ( DownstreamStackBusLane[31][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane22_strm1_data          ( DownstreamStackBusLane[31][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane22_strm1_data_valid    ( DownstreamStackBusLane[31][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane23_strm0_ready         ( DownstreamStackBusLane[31][23].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane23_strm0_cntl          ( DownstreamStackBusLane[31][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane23_strm0_data          ( DownstreamStackBusLane[31][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane23_strm0_data_valid    ( DownstreamStackBusLane[31][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane23_strm1_ready         ( DownstreamStackBusLane[31][23].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane23_strm1_cntl          ( DownstreamStackBusLane[31][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane23_strm1_data          ( DownstreamStackBusLane[31][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane23_strm1_data_valid    ( DownstreamStackBusLane[31][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane24_strm0_ready         ( DownstreamStackBusLane[31][24].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane24_strm0_cntl          ( DownstreamStackBusLane[31][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane24_strm0_data          ( DownstreamStackBusLane[31][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane24_strm0_data_valid    ( DownstreamStackBusLane[31][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane24_strm1_ready         ( DownstreamStackBusLane[31][24].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane24_strm1_cntl          ( DownstreamStackBusLane[31][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane24_strm1_data          ( DownstreamStackBusLane[31][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane24_strm1_data_valid    ( DownstreamStackBusLane[31][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane25_strm0_ready         ( DownstreamStackBusLane[31][25].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane25_strm0_cntl          ( DownstreamStackBusLane[31][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane25_strm0_data          ( DownstreamStackBusLane[31][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane25_strm0_data_valid    ( DownstreamStackBusLane[31][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane25_strm1_ready         ( DownstreamStackBusLane[31][25].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane25_strm1_cntl          ( DownstreamStackBusLane[31][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane25_strm1_data          ( DownstreamStackBusLane[31][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane25_strm1_data_valid    ( DownstreamStackBusLane[31][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane26_strm0_ready         ( DownstreamStackBusLane[31][26].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane26_strm0_cntl          ( DownstreamStackBusLane[31][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane26_strm0_data          ( DownstreamStackBusLane[31][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane26_strm0_data_valid    ( DownstreamStackBusLane[31][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane26_strm1_ready         ( DownstreamStackBusLane[31][26].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane26_strm1_cntl          ( DownstreamStackBusLane[31][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane26_strm1_data          ( DownstreamStackBusLane[31][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane26_strm1_data_valid    ( DownstreamStackBusLane[31][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane27_strm0_ready         ( DownstreamStackBusLane[31][27].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane27_strm0_cntl          ( DownstreamStackBusLane[31][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane27_strm0_data          ( DownstreamStackBusLane[31][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane27_strm0_data_valid    ( DownstreamStackBusLane[31][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane27_strm1_ready         ( DownstreamStackBusLane[31][27].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane27_strm1_cntl          ( DownstreamStackBusLane[31][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane27_strm1_data          ( DownstreamStackBusLane[31][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane27_strm1_data_valid    ( DownstreamStackBusLane[31][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane28_strm0_ready         ( DownstreamStackBusLane[31][28].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane28_strm0_cntl          ( DownstreamStackBusLane[31][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane28_strm0_data          ( DownstreamStackBusLane[31][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane28_strm0_data_valid    ( DownstreamStackBusLane[31][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane28_strm1_ready         ( DownstreamStackBusLane[31][28].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane28_strm1_cntl          ( DownstreamStackBusLane[31][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane28_strm1_data          ( DownstreamStackBusLane[31][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane28_strm1_data_valid    ( DownstreamStackBusLane[31][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane29_strm0_ready         ( DownstreamStackBusLane[31][29].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane29_strm0_cntl          ( DownstreamStackBusLane[31][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane29_strm0_data          ( DownstreamStackBusLane[31][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane29_strm0_data_valid    ( DownstreamStackBusLane[31][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane29_strm1_ready         ( DownstreamStackBusLane[31][29].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane29_strm1_cntl          ( DownstreamStackBusLane[31][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane29_strm1_data          ( DownstreamStackBusLane[31][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane29_strm1_data_valid    ( DownstreamStackBusLane[31][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane30_strm0_ready         ( DownstreamStackBusLane[31][30].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane30_strm0_cntl          ( DownstreamStackBusLane[31][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane30_strm0_data          ( DownstreamStackBusLane[31][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane30_strm0_data_valid    ( DownstreamStackBusLane[31][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane30_strm1_ready         ( DownstreamStackBusLane[31][30].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane30_strm1_cntl          ( DownstreamStackBusLane[31][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane30_strm1_data          ( DownstreamStackBusLane[31][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane30_strm1_data_valid    ( DownstreamStackBusLane[31][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 31, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane31_strm0_ready         ( DownstreamStackBusLane[31][31].pe__std__lane_strm0_ready              ),      
        .std__pe31__lane31_strm0_cntl          ( DownstreamStackBusLane[31][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe31__lane31_strm0_data          ( DownstreamStackBusLane[31][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe31__lane31_strm0_data_valid    ( DownstreamStackBusLane[31][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__std__lane31_strm1_ready         ( DownstreamStackBusLane[31][31].pe__std__lane_strm1_ready              ),      
        .std__pe31__lane31_strm1_cntl          ( DownstreamStackBusLane[31][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe31__lane31_strm1_data          ( DownstreamStackBusLane[31][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe31__lane31_strm1_data_valid    ( DownstreamStackBusLane[31][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane0_strm0_ready         ( DownstreamStackBusLane[32][0].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane0_strm0_cntl          ( DownstreamStackBusLane[32][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane0_strm0_data          ( DownstreamStackBusLane[32][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane0_strm0_data_valid    ( DownstreamStackBusLane[32][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane0_strm1_ready         ( DownstreamStackBusLane[32][0].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane0_strm1_cntl          ( DownstreamStackBusLane[32][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane0_strm1_data          ( DownstreamStackBusLane[32][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane0_strm1_data_valid    ( DownstreamStackBusLane[32][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane1_strm0_ready         ( DownstreamStackBusLane[32][1].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane1_strm0_cntl          ( DownstreamStackBusLane[32][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane1_strm0_data          ( DownstreamStackBusLane[32][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane1_strm0_data_valid    ( DownstreamStackBusLane[32][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane1_strm1_ready         ( DownstreamStackBusLane[32][1].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane1_strm1_cntl          ( DownstreamStackBusLane[32][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane1_strm1_data          ( DownstreamStackBusLane[32][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane1_strm1_data_valid    ( DownstreamStackBusLane[32][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane2_strm0_ready         ( DownstreamStackBusLane[32][2].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane2_strm0_cntl          ( DownstreamStackBusLane[32][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane2_strm0_data          ( DownstreamStackBusLane[32][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane2_strm0_data_valid    ( DownstreamStackBusLane[32][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane2_strm1_ready         ( DownstreamStackBusLane[32][2].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane2_strm1_cntl          ( DownstreamStackBusLane[32][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane2_strm1_data          ( DownstreamStackBusLane[32][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane2_strm1_data_valid    ( DownstreamStackBusLane[32][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane3_strm0_ready         ( DownstreamStackBusLane[32][3].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane3_strm0_cntl          ( DownstreamStackBusLane[32][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane3_strm0_data          ( DownstreamStackBusLane[32][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane3_strm0_data_valid    ( DownstreamStackBusLane[32][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane3_strm1_ready         ( DownstreamStackBusLane[32][3].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane3_strm1_cntl          ( DownstreamStackBusLane[32][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane3_strm1_data          ( DownstreamStackBusLane[32][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane3_strm1_data_valid    ( DownstreamStackBusLane[32][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane4_strm0_ready         ( DownstreamStackBusLane[32][4].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane4_strm0_cntl          ( DownstreamStackBusLane[32][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane4_strm0_data          ( DownstreamStackBusLane[32][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane4_strm0_data_valid    ( DownstreamStackBusLane[32][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane4_strm1_ready         ( DownstreamStackBusLane[32][4].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane4_strm1_cntl          ( DownstreamStackBusLane[32][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane4_strm1_data          ( DownstreamStackBusLane[32][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane4_strm1_data_valid    ( DownstreamStackBusLane[32][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane5_strm0_ready         ( DownstreamStackBusLane[32][5].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane5_strm0_cntl          ( DownstreamStackBusLane[32][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane5_strm0_data          ( DownstreamStackBusLane[32][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane5_strm0_data_valid    ( DownstreamStackBusLane[32][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane5_strm1_ready         ( DownstreamStackBusLane[32][5].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane5_strm1_cntl          ( DownstreamStackBusLane[32][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane5_strm1_data          ( DownstreamStackBusLane[32][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane5_strm1_data_valid    ( DownstreamStackBusLane[32][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane6_strm0_ready         ( DownstreamStackBusLane[32][6].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane6_strm0_cntl          ( DownstreamStackBusLane[32][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane6_strm0_data          ( DownstreamStackBusLane[32][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane6_strm0_data_valid    ( DownstreamStackBusLane[32][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane6_strm1_ready         ( DownstreamStackBusLane[32][6].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane6_strm1_cntl          ( DownstreamStackBusLane[32][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane6_strm1_data          ( DownstreamStackBusLane[32][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane6_strm1_data_valid    ( DownstreamStackBusLane[32][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane7_strm0_ready         ( DownstreamStackBusLane[32][7].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane7_strm0_cntl          ( DownstreamStackBusLane[32][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane7_strm0_data          ( DownstreamStackBusLane[32][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane7_strm0_data_valid    ( DownstreamStackBusLane[32][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane7_strm1_ready         ( DownstreamStackBusLane[32][7].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane7_strm1_cntl          ( DownstreamStackBusLane[32][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane7_strm1_data          ( DownstreamStackBusLane[32][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane7_strm1_data_valid    ( DownstreamStackBusLane[32][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane8_strm0_ready         ( DownstreamStackBusLane[32][8].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane8_strm0_cntl          ( DownstreamStackBusLane[32][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane8_strm0_data          ( DownstreamStackBusLane[32][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane8_strm0_data_valid    ( DownstreamStackBusLane[32][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane8_strm1_ready         ( DownstreamStackBusLane[32][8].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane8_strm1_cntl          ( DownstreamStackBusLane[32][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane8_strm1_data          ( DownstreamStackBusLane[32][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane8_strm1_data_valid    ( DownstreamStackBusLane[32][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane9_strm0_ready         ( DownstreamStackBusLane[32][9].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane9_strm0_cntl          ( DownstreamStackBusLane[32][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane9_strm0_data          ( DownstreamStackBusLane[32][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane9_strm0_data_valid    ( DownstreamStackBusLane[32][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane9_strm1_ready         ( DownstreamStackBusLane[32][9].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane9_strm1_cntl          ( DownstreamStackBusLane[32][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane9_strm1_data          ( DownstreamStackBusLane[32][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane9_strm1_data_valid    ( DownstreamStackBusLane[32][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane10_strm0_ready         ( DownstreamStackBusLane[32][10].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane10_strm0_cntl          ( DownstreamStackBusLane[32][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane10_strm0_data          ( DownstreamStackBusLane[32][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane10_strm0_data_valid    ( DownstreamStackBusLane[32][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane10_strm1_ready         ( DownstreamStackBusLane[32][10].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane10_strm1_cntl          ( DownstreamStackBusLane[32][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane10_strm1_data          ( DownstreamStackBusLane[32][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane10_strm1_data_valid    ( DownstreamStackBusLane[32][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane11_strm0_ready         ( DownstreamStackBusLane[32][11].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane11_strm0_cntl          ( DownstreamStackBusLane[32][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane11_strm0_data          ( DownstreamStackBusLane[32][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane11_strm0_data_valid    ( DownstreamStackBusLane[32][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane11_strm1_ready         ( DownstreamStackBusLane[32][11].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane11_strm1_cntl          ( DownstreamStackBusLane[32][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane11_strm1_data          ( DownstreamStackBusLane[32][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane11_strm1_data_valid    ( DownstreamStackBusLane[32][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane12_strm0_ready         ( DownstreamStackBusLane[32][12].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane12_strm0_cntl          ( DownstreamStackBusLane[32][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane12_strm0_data          ( DownstreamStackBusLane[32][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane12_strm0_data_valid    ( DownstreamStackBusLane[32][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane12_strm1_ready         ( DownstreamStackBusLane[32][12].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane12_strm1_cntl          ( DownstreamStackBusLane[32][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane12_strm1_data          ( DownstreamStackBusLane[32][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane12_strm1_data_valid    ( DownstreamStackBusLane[32][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane13_strm0_ready         ( DownstreamStackBusLane[32][13].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane13_strm0_cntl          ( DownstreamStackBusLane[32][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane13_strm0_data          ( DownstreamStackBusLane[32][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane13_strm0_data_valid    ( DownstreamStackBusLane[32][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane13_strm1_ready         ( DownstreamStackBusLane[32][13].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane13_strm1_cntl          ( DownstreamStackBusLane[32][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane13_strm1_data          ( DownstreamStackBusLane[32][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane13_strm1_data_valid    ( DownstreamStackBusLane[32][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane14_strm0_ready         ( DownstreamStackBusLane[32][14].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane14_strm0_cntl          ( DownstreamStackBusLane[32][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane14_strm0_data          ( DownstreamStackBusLane[32][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane14_strm0_data_valid    ( DownstreamStackBusLane[32][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane14_strm1_ready         ( DownstreamStackBusLane[32][14].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane14_strm1_cntl          ( DownstreamStackBusLane[32][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane14_strm1_data          ( DownstreamStackBusLane[32][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane14_strm1_data_valid    ( DownstreamStackBusLane[32][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane15_strm0_ready         ( DownstreamStackBusLane[32][15].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane15_strm0_cntl          ( DownstreamStackBusLane[32][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane15_strm0_data          ( DownstreamStackBusLane[32][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane15_strm0_data_valid    ( DownstreamStackBusLane[32][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane15_strm1_ready         ( DownstreamStackBusLane[32][15].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane15_strm1_cntl          ( DownstreamStackBusLane[32][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane15_strm1_data          ( DownstreamStackBusLane[32][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane15_strm1_data_valid    ( DownstreamStackBusLane[32][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane16_strm0_ready         ( DownstreamStackBusLane[32][16].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane16_strm0_cntl          ( DownstreamStackBusLane[32][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane16_strm0_data          ( DownstreamStackBusLane[32][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane16_strm0_data_valid    ( DownstreamStackBusLane[32][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane16_strm1_ready         ( DownstreamStackBusLane[32][16].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane16_strm1_cntl          ( DownstreamStackBusLane[32][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane16_strm1_data          ( DownstreamStackBusLane[32][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane16_strm1_data_valid    ( DownstreamStackBusLane[32][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane17_strm0_ready         ( DownstreamStackBusLane[32][17].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane17_strm0_cntl          ( DownstreamStackBusLane[32][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane17_strm0_data          ( DownstreamStackBusLane[32][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane17_strm0_data_valid    ( DownstreamStackBusLane[32][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane17_strm1_ready         ( DownstreamStackBusLane[32][17].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane17_strm1_cntl          ( DownstreamStackBusLane[32][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane17_strm1_data          ( DownstreamStackBusLane[32][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane17_strm1_data_valid    ( DownstreamStackBusLane[32][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane18_strm0_ready         ( DownstreamStackBusLane[32][18].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane18_strm0_cntl          ( DownstreamStackBusLane[32][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane18_strm0_data          ( DownstreamStackBusLane[32][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane18_strm0_data_valid    ( DownstreamStackBusLane[32][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane18_strm1_ready         ( DownstreamStackBusLane[32][18].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane18_strm1_cntl          ( DownstreamStackBusLane[32][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane18_strm1_data          ( DownstreamStackBusLane[32][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane18_strm1_data_valid    ( DownstreamStackBusLane[32][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane19_strm0_ready         ( DownstreamStackBusLane[32][19].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane19_strm0_cntl          ( DownstreamStackBusLane[32][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane19_strm0_data          ( DownstreamStackBusLane[32][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane19_strm0_data_valid    ( DownstreamStackBusLane[32][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane19_strm1_ready         ( DownstreamStackBusLane[32][19].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane19_strm1_cntl          ( DownstreamStackBusLane[32][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane19_strm1_data          ( DownstreamStackBusLane[32][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane19_strm1_data_valid    ( DownstreamStackBusLane[32][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane20_strm0_ready         ( DownstreamStackBusLane[32][20].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane20_strm0_cntl          ( DownstreamStackBusLane[32][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane20_strm0_data          ( DownstreamStackBusLane[32][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane20_strm0_data_valid    ( DownstreamStackBusLane[32][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane20_strm1_ready         ( DownstreamStackBusLane[32][20].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane20_strm1_cntl          ( DownstreamStackBusLane[32][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane20_strm1_data          ( DownstreamStackBusLane[32][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane20_strm1_data_valid    ( DownstreamStackBusLane[32][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane21_strm0_ready         ( DownstreamStackBusLane[32][21].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane21_strm0_cntl          ( DownstreamStackBusLane[32][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane21_strm0_data          ( DownstreamStackBusLane[32][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane21_strm0_data_valid    ( DownstreamStackBusLane[32][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane21_strm1_ready         ( DownstreamStackBusLane[32][21].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane21_strm1_cntl          ( DownstreamStackBusLane[32][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane21_strm1_data          ( DownstreamStackBusLane[32][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane21_strm1_data_valid    ( DownstreamStackBusLane[32][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane22_strm0_ready         ( DownstreamStackBusLane[32][22].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane22_strm0_cntl          ( DownstreamStackBusLane[32][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane22_strm0_data          ( DownstreamStackBusLane[32][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane22_strm0_data_valid    ( DownstreamStackBusLane[32][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane22_strm1_ready         ( DownstreamStackBusLane[32][22].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane22_strm1_cntl          ( DownstreamStackBusLane[32][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane22_strm1_data          ( DownstreamStackBusLane[32][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane22_strm1_data_valid    ( DownstreamStackBusLane[32][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane23_strm0_ready         ( DownstreamStackBusLane[32][23].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane23_strm0_cntl          ( DownstreamStackBusLane[32][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane23_strm0_data          ( DownstreamStackBusLane[32][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane23_strm0_data_valid    ( DownstreamStackBusLane[32][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane23_strm1_ready         ( DownstreamStackBusLane[32][23].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane23_strm1_cntl          ( DownstreamStackBusLane[32][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane23_strm1_data          ( DownstreamStackBusLane[32][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane23_strm1_data_valid    ( DownstreamStackBusLane[32][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane24_strm0_ready         ( DownstreamStackBusLane[32][24].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane24_strm0_cntl          ( DownstreamStackBusLane[32][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane24_strm0_data          ( DownstreamStackBusLane[32][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane24_strm0_data_valid    ( DownstreamStackBusLane[32][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane24_strm1_ready         ( DownstreamStackBusLane[32][24].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane24_strm1_cntl          ( DownstreamStackBusLane[32][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane24_strm1_data          ( DownstreamStackBusLane[32][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane24_strm1_data_valid    ( DownstreamStackBusLane[32][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane25_strm0_ready         ( DownstreamStackBusLane[32][25].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane25_strm0_cntl          ( DownstreamStackBusLane[32][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane25_strm0_data          ( DownstreamStackBusLane[32][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane25_strm0_data_valid    ( DownstreamStackBusLane[32][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane25_strm1_ready         ( DownstreamStackBusLane[32][25].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane25_strm1_cntl          ( DownstreamStackBusLane[32][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane25_strm1_data          ( DownstreamStackBusLane[32][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane25_strm1_data_valid    ( DownstreamStackBusLane[32][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane26_strm0_ready         ( DownstreamStackBusLane[32][26].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane26_strm0_cntl          ( DownstreamStackBusLane[32][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane26_strm0_data          ( DownstreamStackBusLane[32][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane26_strm0_data_valid    ( DownstreamStackBusLane[32][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane26_strm1_ready         ( DownstreamStackBusLane[32][26].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane26_strm1_cntl          ( DownstreamStackBusLane[32][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane26_strm1_data          ( DownstreamStackBusLane[32][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane26_strm1_data_valid    ( DownstreamStackBusLane[32][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane27_strm0_ready         ( DownstreamStackBusLane[32][27].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane27_strm0_cntl          ( DownstreamStackBusLane[32][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane27_strm0_data          ( DownstreamStackBusLane[32][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane27_strm0_data_valid    ( DownstreamStackBusLane[32][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane27_strm1_ready         ( DownstreamStackBusLane[32][27].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane27_strm1_cntl          ( DownstreamStackBusLane[32][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane27_strm1_data          ( DownstreamStackBusLane[32][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane27_strm1_data_valid    ( DownstreamStackBusLane[32][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane28_strm0_ready         ( DownstreamStackBusLane[32][28].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane28_strm0_cntl          ( DownstreamStackBusLane[32][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane28_strm0_data          ( DownstreamStackBusLane[32][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane28_strm0_data_valid    ( DownstreamStackBusLane[32][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane28_strm1_ready         ( DownstreamStackBusLane[32][28].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane28_strm1_cntl          ( DownstreamStackBusLane[32][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane28_strm1_data          ( DownstreamStackBusLane[32][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane28_strm1_data_valid    ( DownstreamStackBusLane[32][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane29_strm0_ready         ( DownstreamStackBusLane[32][29].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane29_strm0_cntl          ( DownstreamStackBusLane[32][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane29_strm0_data          ( DownstreamStackBusLane[32][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane29_strm0_data_valid    ( DownstreamStackBusLane[32][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane29_strm1_ready         ( DownstreamStackBusLane[32][29].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane29_strm1_cntl          ( DownstreamStackBusLane[32][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane29_strm1_data          ( DownstreamStackBusLane[32][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane29_strm1_data_valid    ( DownstreamStackBusLane[32][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane30_strm0_ready         ( DownstreamStackBusLane[32][30].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane30_strm0_cntl          ( DownstreamStackBusLane[32][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane30_strm0_data          ( DownstreamStackBusLane[32][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane30_strm0_data_valid    ( DownstreamStackBusLane[32][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane30_strm1_ready         ( DownstreamStackBusLane[32][30].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane30_strm1_cntl          ( DownstreamStackBusLane[32][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane30_strm1_data          ( DownstreamStackBusLane[32][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane30_strm1_data_valid    ( DownstreamStackBusLane[32][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 32, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane31_strm0_ready         ( DownstreamStackBusLane[32][31].pe__std__lane_strm0_ready              ),      
        .std__pe32__lane31_strm0_cntl          ( DownstreamStackBusLane[32][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe32__lane31_strm0_data          ( DownstreamStackBusLane[32][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe32__lane31_strm0_data_valid    ( DownstreamStackBusLane[32][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__std__lane31_strm1_ready         ( DownstreamStackBusLane[32][31].pe__std__lane_strm1_ready              ),      
        .std__pe32__lane31_strm1_cntl          ( DownstreamStackBusLane[32][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe32__lane31_strm1_data          ( DownstreamStackBusLane[32][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe32__lane31_strm1_data_valid    ( DownstreamStackBusLane[32][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane0_strm0_ready         ( DownstreamStackBusLane[33][0].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane0_strm0_cntl          ( DownstreamStackBusLane[33][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane0_strm0_data          ( DownstreamStackBusLane[33][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane0_strm0_data_valid    ( DownstreamStackBusLane[33][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane0_strm1_ready         ( DownstreamStackBusLane[33][0].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane0_strm1_cntl          ( DownstreamStackBusLane[33][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane0_strm1_data          ( DownstreamStackBusLane[33][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane0_strm1_data_valid    ( DownstreamStackBusLane[33][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane1_strm0_ready         ( DownstreamStackBusLane[33][1].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane1_strm0_cntl          ( DownstreamStackBusLane[33][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane1_strm0_data          ( DownstreamStackBusLane[33][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane1_strm0_data_valid    ( DownstreamStackBusLane[33][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane1_strm1_ready         ( DownstreamStackBusLane[33][1].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane1_strm1_cntl          ( DownstreamStackBusLane[33][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane1_strm1_data          ( DownstreamStackBusLane[33][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane1_strm1_data_valid    ( DownstreamStackBusLane[33][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane2_strm0_ready         ( DownstreamStackBusLane[33][2].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane2_strm0_cntl          ( DownstreamStackBusLane[33][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane2_strm0_data          ( DownstreamStackBusLane[33][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane2_strm0_data_valid    ( DownstreamStackBusLane[33][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane2_strm1_ready         ( DownstreamStackBusLane[33][2].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane2_strm1_cntl          ( DownstreamStackBusLane[33][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane2_strm1_data          ( DownstreamStackBusLane[33][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane2_strm1_data_valid    ( DownstreamStackBusLane[33][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane3_strm0_ready         ( DownstreamStackBusLane[33][3].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane3_strm0_cntl          ( DownstreamStackBusLane[33][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane3_strm0_data          ( DownstreamStackBusLane[33][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane3_strm0_data_valid    ( DownstreamStackBusLane[33][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane3_strm1_ready         ( DownstreamStackBusLane[33][3].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane3_strm1_cntl          ( DownstreamStackBusLane[33][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane3_strm1_data          ( DownstreamStackBusLane[33][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane3_strm1_data_valid    ( DownstreamStackBusLane[33][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane4_strm0_ready         ( DownstreamStackBusLane[33][4].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane4_strm0_cntl          ( DownstreamStackBusLane[33][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane4_strm0_data          ( DownstreamStackBusLane[33][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane4_strm0_data_valid    ( DownstreamStackBusLane[33][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane4_strm1_ready         ( DownstreamStackBusLane[33][4].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane4_strm1_cntl          ( DownstreamStackBusLane[33][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane4_strm1_data          ( DownstreamStackBusLane[33][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane4_strm1_data_valid    ( DownstreamStackBusLane[33][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane5_strm0_ready         ( DownstreamStackBusLane[33][5].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane5_strm0_cntl          ( DownstreamStackBusLane[33][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane5_strm0_data          ( DownstreamStackBusLane[33][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane5_strm0_data_valid    ( DownstreamStackBusLane[33][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane5_strm1_ready         ( DownstreamStackBusLane[33][5].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane5_strm1_cntl          ( DownstreamStackBusLane[33][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane5_strm1_data          ( DownstreamStackBusLane[33][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane5_strm1_data_valid    ( DownstreamStackBusLane[33][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane6_strm0_ready         ( DownstreamStackBusLane[33][6].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane6_strm0_cntl          ( DownstreamStackBusLane[33][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane6_strm0_data          ( DownstreamStackBusLane[33][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane6_strm0_data_valid    ( DownstreamStackBusLane[33][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane6_strm1_ready         ( DownstreamStackBusLane[33][6].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane6_strm1_cntl          ( DownstreamStackBusLane[33][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane6_strm1_data          ( DownstreamStackBusLane[33][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane6_strm1_data_valid    ( DownstreamStackBusLane[33][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane7_strm0_ready         ( DownstreamStackBusLane[33][7].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane7_strm0_cntl          ( DownstreamStackBusLane[33][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane7_strm0_data          ( DownstreamStackBusLane[33][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane7_strm0_data_valid    ( DownstreamStackBusLane[33][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane7_strm1_ready         ( DownstreamStackBusLane[33][7].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane7_strm1_cntl          ( DownstreamStackBusLane[33][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane7_strm1_data          ( DownstreamStackBusLane[33][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane7_strm1_data_valid    ( DownstreamStackBusLane[33][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane8_strm0_ready         ( DownstreamStackBusLane[33][8].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane8_strm0_cntl          ( DownstreamStackBusLane[33][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane8_strm0_data          ( DownstreamStackBusLane[33][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane8_strm0_data_valid    ( DownstreamStackBusLane[33][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane8_strm1_ready         ( DownstreamStackBusLane[33][8].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane8_strm1_cntl          ( DownstreamStackBusLane[33][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane8_strm1_data          ( DownstreamStackBusLane[33][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane8_strm1_data_valid    ( DownstreamStackBusLane[33][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane9_strm0_ready         ( DownstreamStackBusLane[33][9].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane9_strm0_cntl          ( DownstreamStackBusLane[33][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane9_strm0_data          ( DownstreamStackBusLane[33][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane9_strm0_data_valid    ( DownstreamStackBusLane[33][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane9_strm1_ready         ( DownstreamStackBusLane[33][9].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane9_strm1_cntl          ( DownstreamStackBusLane[33][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane9_strm1_data          ( DownstreamStackBusLane[33][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane9_strm1_data_valid    ( DownstreamStackBusLane[33][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane10_strm0_ready         ( DownstreamStackBusLane[33][10].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane10_strm0_cntl          ( DownstreamStackBusLane[33][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane10_strm0_data          ( DownstreamStackBusLane[33][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane10_strm0_data_valid    ( DownstreamStackBusLane[33][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane10_strm1_ready         ( DownstreamStackBusLane[33][10].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane10_strm1_cntl          ( DownstreamStackBusLane[33][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane10_strm1_data          ( DownstreamStackBusLane[33][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane10_strm1_data_valid    ( DownstreamStackBusLane[33][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane11_strm0_ready         ( DownstreamStackBusLane[33][11].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane11_strm0_cntl          ( DownstreamStackBusLane[33][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane11_strm0_data          ( DownstreamStackBusLane[33][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane11_strm0_data_valid    ( DownstreamStackBusLane[33][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane11_strm1_ready         ( DownstreamStackBusLane[33][11].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane11_strm1_cntl          ( DownstreamStackBusLane[33][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane11_strm1_data          ( DownstreamStackBusLane[33][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane11_strm1_data_valid    ( DownstreamStackBusLane[33][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane12_strm0_ready         ( DownstreamStackBusLane[33][12].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane12_strm0_cntl          ( DownstreamStackBusLane[33][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane12_strm0_data          ( DownstreamStackBusLane[33][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane12_strm0_data_valid    ( DownstreamStackBusLane[33][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane12_strm1_ready         ( DownstreamStackBusLane[33][12].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane12_strm1_cntl          ( DownstreamStackBusLane[33][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane12_strm1_data          ( DownstreamStackBusLane[33][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane12_strm1_data_valid    ( DownstreamStackBusLane[33][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane13_strm0_ready         ( DownstreamStackBusLane[33][13].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane13_strm0_cntl          ( DownstreamStackBusLane[33][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane13_strm0_data          ( DownstreamStackBusLane[33][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane13_strm0_data_valid    ( DownstreamStackBusLane[33][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane13_strm1_ready         ( DownstreamStackBusLane[33][13].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane13_strm1_cntl          ( DownstreamStackBusLane[33][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane13_strm1_data          ( DownstreamStackBusLane[33][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane13_strm1_data_valid    ( DownstreamStackBusLane[33][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane14_strm0_ready         ( DownstreamStackBusLane[33][14].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane14_strm0_cntl          ( DownstreamStackBusLane[33][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane14_strm0_data          ( DownstreamStackBusLane[33][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane14_strm0_data_valid    ( DownstreamStackBusLane[33][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane14_strm1_ready         ( DownstreamStackBusLane[33][14].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane14_strm1_cntl          ( DownstreamStackBusLane[33][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane14_strm1_data          ( DownstreamStackBusLane[33][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane14_strm1_data_valid    ( DownstreamStackBusLane[33][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane15_strm0_ready         ( DownstreamStackBusLane[33][15].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane15_strm0_cntl          ( DownstreamStackBusLane[33][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane15_strm0_data          ( DownstreamStackBusLane[33][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane15_strm0_data_valid    ( DownstreamStackBusLane[33][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane15_strm1_ready         ( DownstreamStackBusLane[33][15].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane15_strm1_cntl          ( DownstreamStackBusLane[33][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane15_strm1_data          ( DownstreamStackBusLane[33][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane15_strm1_data_valid    ( DownstreamStackBusLane[33][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane16_strm0_ready         ( DownstreamStackBusLane[33][16].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane16_strm0_cntl          ( DownstreamStackBusLane[33][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane16_strm0_data          ( DownstreamStackBusLane[33][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane16_strm0_data_valid    ( DownstreamStackBusLane[33][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane16_strm1_ready         ( DownstreamStackBusLane[33][16].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane16_strm1_cntl          ( DownstreamStackBusLane[33][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane16_strm1_data          ( DownstreamStackBusLane[33][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane16_strm1_data_valid    ( DownstreamStackBusLane[33][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane17_strm0_ready         ( DownstreamStackBusLane[33][17].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane17_strm0_cntl          ( DownstreamStackBusLane[33][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane17_strm0_data          ( DownstreamStackBusLane[33][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane17_strm0_data_valid    ( DownstreamStackBusLane[33][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane17_strm1_ready         ( DownstreamStackBusLane[33][17].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane17_strm1_cntl          ( DownstreamStackBusLane[33][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane17_strm1_data          ( DownstreamStackBusLane[33][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane17_strm1_data_valid    ( DownstreamStackBusLane[33][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane18_strm0_ready         ( DownstreamStackBusLane[33][18].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane18_strm0_cntl          ( DownstreamStackBusLane[33][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane18_strm0_data          ( DownstreamStackBusLane[33][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane18_strm0_data_valid    ( DownstreamStackBusLane[33][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane18_strm1_ready         ( DownstreamStackBusLane[33][18].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane18_strm1_cntl          ( DownstreamStackBusLane[33][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane18_strm1_data          ( DownstreamStackBusLane[33][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane18_strm1_data_valid    ( DownstreamStackBusLane[33][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane19_strm0_ready         ( DownstreamStackBusLane[33][19].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane19_strm0_cntl          ( DownstreamStackBusLane[33][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane19_strm0_data          ( DownstreamStackBusLane[33][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane19_strm0_data_valid    ( DownstreamStackBusLane[33][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane19_strm1_ready         ( DownstreamStackBusLane[33][19].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane19_strm1_cntl          ( DownstreamStackBusLane[33][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane19_strm1_data          ( DownstreamStackBusLane[33][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane19_strm1_data_valid    ( DownstreamStackBusLane[33][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane20_strm0_ready         ( DownstreamStackBusLane[33][20].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane20_strm0_cntl          ( DownstreamStackBusLane[33][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane20_strm0_data          ( DownstreamStackBusLane[33][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane20_strm0_data_valid    ( DownstreamStackBusLane[33][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane20_strm1_ready         ( DownstreamStackBusLane[33][20].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane20_strm1_cntl          ( DownstreamStackBusLane[33][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane20_strm1_data          ( DownstreamStackBusLane[33][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane20_strm1_data_valid    ( DownstreamStackBusLane[33][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane21_strm0_ready         ( DownstreamStackBusLane[33][21].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane21_strm0_cntl          ( DownstreamStackBusLane[33][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane21_strm0_data          ( DownstreamStackBusLane[33][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane21_strm0_data_valid    ( DownstreamStackBusLane[33][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane21_strm1_ready         ( DownstreamStackBusLane[33][21].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane21_strm1_cntl          ( DownstreamStackBusLane[33][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane21_strm1_data          ( DownstreamStackBusLane[33][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane21_strm1_data_valid    ( DownstreamStackBusLane[33][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane22_strm0_ready         ( DownstreamStackBusLane[33][22].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane22_strm0_cntl          ( DownstreamStackBusLane[33][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane22_strm0_data          ( DownstreamStackBusLane[33][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane22_strm0_data_valid    ( DownstreamStackBusLane[33][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane22_strm1_ready         ( DownstreamStackBusLane[33][22].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane22_strm1_cntl          ( DownstreamStackBusLane[33][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane22_strm1_data          ( DownstreamStackBusLane[33][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane22_strm1_data_valid    ( DownstreamStackBusLane[33][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane23_strm0_ready         ( DownstreamStackBusLane[33][23].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane23_strm0_cntl          ( DownstreamStackBusLane[33][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane23_strm0_data          ( DownstreamStackBusLane[33][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane23_strm0_data_valid    ( DownstreamStackBusLane[33][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane23_strm1_ready         ( DownstreamStackBusLane[33][23].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane23_strm1_cntl          ( DownstreamStackBusLane[33][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane23_strm1_data          ( DownstreamStackBusLane[33][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane23_strm1_data_valid    ( DownstreamStackBusLane[33][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane24_strm0_ready         ( DownstreamStackBusLane[33][24].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane24_strm0_cntl          ( DownstreamStackBusLane[33][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane24_strm0_data          ( DownstreamStackBusLane[33][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane24_strm0_data_valid    ( DownstreamStackBusLane[33][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane24_strm1_ready         ( DownstreamStackBusLane[33][24].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane24_strm1_cntl          ( DownstreamStackBusLane[33][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane24_strm1_data          ( DownstreamStackBusLane[33][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane24_strm1_data_valid    ( DownstreamStackBusLane[33][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane25_strm0_ready         ( DownstreamStackBusLane[33][25].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane25_strm0_cntl          ( DownstreamStackBusLane[33][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane25_strm0_data          ( DownstreamStackBusLane[33][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane25_strm0_data_valid    ( DownstreamStackBusLane[33][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane25_strm1_ready         ( DownstreamStackBusLane[33][25].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane25_strm1_cntl          ( DownstreamStackBusLane[33][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane25_strm1_data          ( DownstreamStackBusLane[33][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane25_strm1_data_valid    ( DownstreamStackBusLane[33][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane26_strm0_ready         ( DownstreamStackBusLane[33][26].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane26_strm0_cntl          ( DownstreamStackBusLane[33][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane26_strm0_data          ( DownstreamStackBusLane[33][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane26_strm0_data_valid    ( DownstreamStackBusLane[33][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane26_strm1_ready         ( DownstreamStackBusLane[33][26].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane26_strm1_cntl          ( DownstreamStackBusLane[33][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane26_strm1_data          ( DownstreamStackBusLane[33][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane26_strm1_data_valid    ( DownstreamStackBusLane[33][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane27_strm0_ready         ( DownstreamStackBusLane[33][27].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane27_strm0_cntl          ( DownstreamStackBusLane[33][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane27_strm0_data          ( DownstreamStackBusLane[33][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane27_strm0_data_valid    ( DownstreamStackBusLane[33][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane27_strm1_ready         ( DownstreamStackBusLane[33][27].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane27_strm1_cntl          ( DownstreamStackBusLane[33][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane27_strm1_data          ( DownstreamStackBusLane[33][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane27_strm1_data_valid    ( DownstreamStackBusLane[33][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane28_strm0_ready         ( DownstreamStackBusLane[33][28].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane28_strm0_cntl          ( DownstreamStackBusLane[33][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane28_strm0_data          ( DownstreamStackBusLane[33][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane28_strm0_data_valid    ( DownstreamStackBusLane[33][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane28_strm1_ready         ( DownstreamStackBusLane[33][28].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane28_strm1_cntl          ( DownstreamStackBusLane[33][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane28_strm1_data          ( DownstreamStackBusLane[33][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane28_strm1_data_valid    ( DownstreamStackBusLane[33][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane29_strm0_ready         ( DownstreamStackBusLane[33][29].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane29_strm0_cntl          ( DownstreamStackBusLane[33][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane29_strm0_data          ( DownstreamStackBusLane[33][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane29_strm0_data_valid    ( DownstreamStackBusLane[33][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane29_strm1_ready         ( DownstreamStackBusLane[33][29].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane29_strm1_cntl          ( DownstreamStackBusLane[33][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane29_strm1_data          ( DownstreamStackBusLane[33][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane29_strm1_data_valid    ( DownstreamStackBusLane[33][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane30_strm0_ready         ( DownstreamStackBusLane[33][30].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane30_strm0_cntl          ( DownstreamStackBusLane[33][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane30_strm0_data          ( DownstreamStackBusLane[33][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane30_strm0_data_valid    ( DownstreamStackBusLane[33][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane30_strm1_ready         ( DownstreamStackBusLane[33][30].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane30_strm1_cntl          ( DownstreamStackBusLane[33][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane30_strm1_data          ( DownstreamStackBusLane[33][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane30_strm1_data_valid    ( DownstreamStackBusLane[33][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 33, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane31_strm0_ready         ( DownstreamStackBusLane[33][31].pe__std__lane_strm0_ready              ),      
        .std__pe33__lane31_strm0_cntl          ( DownstreamStackBusLane[33][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe33__lane31_strm0_data          ( DownstreamStackBusLane[33][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe33__lane31_strm0_data_valid    ( DownstreamStackBusLane[33][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__std__lane31_strm1_ready         ( DownstreamStackBusLane[33][31].pe__std__lane_strm1_ready              ),      
        .std__pe33__lane31_strm1_cntl          ( DownstreamStackBusLane[33][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe33__lane31_strm1_data          ( DownstreamStackBusLane[33][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe33__lane31_strm1_data_valid    ( DownstreamStackBusLane[33][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane0_strm0_ready         ( DownstreamStackBusLane[34][0].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane0_strm0_cntl          ( DownstreamStackBusLane[34][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane0_strm0_data          ( DownstreamStackBusLane[34][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane0_strm0_data_valid    ( DownstreamStackBusLane[34][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane0_strm1_ready         ( DownstreamStackBusLane[34][0].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane0_strm1_cntl          ( DownstreamStackBusLane[34][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane0_strm1_data          ( DownstreamStackBusLane[34][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane0_strm1_data_valid    ( DownstreamStackBusLane[34][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane1_strm0_ready         ( DownstreamStackBusLane[34][1].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane1_strm0_cntl          ( DownstreamStackBusLane[34][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane1_strm0_data          ( DownstreamStackBusLane[34][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane1_strm0_data_valid    ( DownstreamStackBusLane[34][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane1_strm1_ready         ( DownstreamStackBusLane[34][1].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane1_strm1_cntl          ( DownstreamStackBusLane[34][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane1_strm1_data          ( DownstreamStackBusLane[34][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane1_strm1_data_valid    ( DownstreamStackBusLane[34][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane2_strm0_ready         ( DownstreamStackBusLane[34][2].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane2_strm0_cntl          ( DownstreamStackBusLane[34][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane2_strm0_data          ( DownstreamStackBusLane[34][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane2_strm0_data_valid    ( DownstreamStackBusLane[34][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane2_strm1_ready         ( DownstreamStackBusLane[34][2].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane2_strm1_cntl          ( DownstreamStackBusLane[34][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane2_strm1_data          ( DownstreamStackBusLane[34][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane2_strm1_data_valid    ( DownstreamStackBusLane[34][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane3_strm0_ready         ( DownstreamStackBusLane[34][3].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane3_strm0_cntl          ( DownstreamStackBusLane[34][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane3_strm0_data          ( DownstreamStackBusLane[34][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane3_strm0_data_valid    ( DownstreamStackBusLane[34][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane3_strm1_ready         ( DownstreamStackBusLane[34][3].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane3_strm1_cntl          ( DownstreamStackBusLane[34][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane3_strm1_data          ( DownstreamStackBusLane[34][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane3_strm1_data_valid    ( DownstreamStackBusLane[34][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane4_strm0_ready         ( DownstreamStackBusLane[34][4].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane4_strm0_cntl          ( DownstreamStackBusLane[34][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane4_strm0_data          ( DownstreamStackBusLane[34][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane4_strm0_data_valid    ( DownstreamStackBusLane[34][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane4_strm1_ready         ( DownstreamStackBusLane[34][4].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane4_strm1_cntl          ( DownstreamStackBusLane[34][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane4_strm1_data          ( DownstreamStackBusLane[34][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane4_strm1_data_valid    ( DownstreamStackBusLane[34][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane5_strm0_ready         ( DownstreamStackBusLane[34][5].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane5_strm0_cntl          ( DownstreamStackBusLane[34][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane5_strm0_data          ( DownstreamStackBusLane[34][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane5_strm0_data_valid    ( DownstreamStackBusLane[34][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane5_strm1_ready         ( DownstreamStackBusLane[34][5].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane5_strm1_cntl          ( DownstreamStackBusLane[34][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane5_strm1_data          ( DownstreamStackBusLane[34][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane5_strm1_data_valid    ( DownstreamStackBusLane[34][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane6_strm0_ready         ( DownstreamStackBusLane[34][6].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane6_strm0_cntl          ( DownstreamStackBusLane[34][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane6_strm0_data          ( DownstreamStackBusLane[34][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane6_strm0_data_valid    ( DownstreamStackBusLane[34][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane6_strm1_ready         ( DownstreamStackBusLane[34][6].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane6_strm1_cntl          ( DownstreamStackBusLane[34][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane6_strm1_data          ( DownstreamStackBusLane[34][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane6_strm1_data_valid    ( DownstreamStackBusLane[34][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane7_strm0_ready         ( DownstreamStackBusLane[34][7].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane7_strm0_cntl          ( DownstreamStackBusLane[34][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane7_strm0_data          ( DownstreamStackBusLane[34][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane7_strm0_data_valid    ( DownstreamStackBusLane[34][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane7_strm1_ready         ( DownstreamStackBusLane[34][7].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane7_strm1_cntl          ( DownstreamStackBusLane[34][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane7_strm1_data          ( DownstreamStackBusLane[34][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane7_strm1_data_valid    ( DownstreamStackBusLane[34][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane8_strm0_ready         ( DownstreamStackBusLane[34][8].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane8_strm0_cntl          ( DownstreamStackBusLane[34][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane8_strm0_data          ( DownstreamStackBusLane[34][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane8_strm0_data_valid    ( DownstreamStackBusLane[34][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane8_strm1_ready         ( DownstreamStackBusLane[34][8].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane8_strm1_cntl          ( DownstreamStackBusLane[34][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane8_strm1_data          ( DownstreamStackBusLane[34][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane8_strm1_data_valid    ( DownstreamStackBusLane[34][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane9_strm0_ready         ( DownstreamStackBusLane[34][9].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane9_strm0_cntl          ( DownstreamStackBusLane[34][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane9_strm0_data          ( DownstreamStackBusLane[34][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane9_strm0_data_valid    ( DownstreamStackBusLane[34][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane9_strm1_ready         ( DownstreamStackBusLane[34][9].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane9_strm1_cntl          ( DownstreamStackBusLane[34][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane9_strm1_data          ( DownstreamStackBusLane[34][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane9_strm1_data_valid    ( DownstreamStackBusLane[34][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane10_strm0_ready         ( DownstreamStackBusLane[34][10].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane10_strm0_cntl          ( DownstreamStackBusLane[34][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane10_strm0_data          ( DownstreamStackBusLane[34][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane10_strm0_data_valid    ( DownstreamStackBusLane[34][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane10_strm1_ready         ( DownstreamStackBusLane[34][10].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane10_strm1_cntl          ( DownstreamStackBusLane[34][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane10_strm1_data          ( DownstreamStackBusLane[34][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane10_strm1_data_valid    ( DownstreamStackBusLane[34][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane11_strm0_ready         ( DownstreamStackBusLane[34][11].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane11_strm0_cntl          ( DownstreamStackBusLane[34][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane11_strm0_data          ( DownstreamStackBusLane[34][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane11_strm0_data_valid    ( DownstreamStackBusLane[34][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane11_strm1_ready         ( DownstreamStackBusLane[34][11].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane11_strm1_cntl          ( DownstreamStackBusLane[34][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane11_strm1_data          ( DownstreamStackBusLane[34][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane11_strm1_data_valid    ( DownstreamStackBusLane[34][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane12_strm0_ready         ( DownstreamStackBusLane[34][12].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane12_strm0_cntl          ( DownstreamStackBusLane[34][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane12_strm0_data          ( DownstreamStackBusLane[34][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane12_strm0_data_valid    ( DownstreamStackBusLane[34][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane12_strm1_ready         ( DownstreamStackBusLane[34][12].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane12_strm1_cntl          ( DownstreamStackBusLane[34][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane12_strm1_data          ( DownstreamStackBusLane[34][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane12_strm1_data_valid    ( DownstreamStackBusLane[34][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane13_strm0_ready         ( DownstreamStackBusLane[34][13].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane13_strm0_cntl          ( DownstreamStackBusLane[34][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane13_strm0_data          ( DownstreamStackBusLane[34][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane13_strm0_data_valid    ( DownstreamStackBusLane[34][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane13_strm1_ready         ( DownstreamStackBusLane[34][13].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane13_strm1_cntl          ( DownstreamStackBusLane[34][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane13_strm1_data          ( DownstreamStackBusLane[34][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane13_strm1_data_valid    ( DownstreamStackBusLane[34][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane14_strm0_ready         ( DownstreamStackBusLane[34][14].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane14_strm0_cntl          ( DownstreamStackBusLane[34][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane14_strm0_data          ( DownstreamStackBusLane[34][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane14_strm0_data_valid    ( DownstreamStackBusLane[34][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane14_strm1_ready         ( DownstreamStackBusLane[34][14].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane14_strm1_cntl          ( DownstreamStackBusLane[34][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane14_strm1_data          ( DownstreamStackBusLane[34][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane14_strm1_data_valid    ( DownstreamStackBusLane[34][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane15_strm0_ready         ( DownstreamStackBusLane[34][15].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane15_strm0_cntl          ( DownstreamStackBusLane[34][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane15_strm0_data          ( DownstreamStackBusLane[34][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane15_strm0_data_valid    ( DownstreamStackBusLane[34][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane15_strm1_ready         ( DownstreamStackBusLane[34][15].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane15_strm1_cntl          ( DownstreamStackBusLane[34][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane15_strm1_data          ( DownstreamStackBusLane[34][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane15_strm1_data_valid    ( DownstreamStackBusLane[34][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane16_strm0_ready         ( DownstreamStackBusLane[34][16].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane16_strm0_cntl          ( DownstreamStackBusLane[34][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane16_strm0_data          ( DownstreamStackBusLane[34][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane16_strm0_data_valid    ( DownstreamStackBusLane[34][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane16_strm1_ready         ( DownstreamStackBusLane[34][16].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane16_strm1_cntl          ( DownstreamStackBusLane[34][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane16_strm1_data          ( DownstreamStackBusLane[34][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane16_strm1_data_valid    ( DownstreamStackBusLane[34][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane17_strm0_ready         ( DownstreamStackBusLane[34][17].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane17_strm0_cntl          ( DownstreamStackBusLane[34][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane17_strm0_data          ( DownstreamStackBusLane[34][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane17_strm0_data_valid    ( DownstreamStackBusLane[34][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane17_strm1_ready         ( DownstreamStackBusLane[34][17].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane17_strm1_cntl          ( DownstreamStackBusLane[34][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane17_strm1_data          ( DownstreamStackBusLane[34][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane17_strm1_data_valid    ( DownstreamStackBusLane[34][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane18_strm0_ready         ( DownstreamStackBusLane[34][18].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane18_strm0_cntl          ( DownstreamStackBusLane[34][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane18_strm0_data          ( DownstreamStackBusLane[34][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane18_strm0_data_valid    ( DownstreamStackBusLane[34][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane18_strm1_ready         ( DownstreamStackBusLane[34][18].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane18_strm1_cntl          ( DownstreamStackBusLane[34][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane18_strm1_data          ( DownstreamStackBusLane[34][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane18_strm1_data_valid    ( DownstreamStackBusLane[34][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane19_strm0_ready         ( DownstreamStackBusLane[34][19].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane19_strm0_cntl          ( DownstreamStackBusLane[34][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane19_strm0_data          ( DownstreamStackBusLane[34][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane19_strm0_data_valid    ( DownstreamStackBusLane[34][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane19_strm1_ready         ( DownstreamStackBusLane[34][19].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane19_strm1_cntl          ( DownstreamStackBusLane[34][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane19_strm1_data          ( DownstreamStackBusLane[34][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane19_strm1_data_valid    ( DownstreamStackBusLane[34][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane20_strm0_ready         ( DownstreamStackBusLane[34][20].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane20_strm0_cntl          ( DownstreamStackBusLane[34][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane20_strm0_data          ( DownstreamStackBusLane[34][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane20_strm0_data_valid    ( DownstreamStackBusLane[34][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane20_strm1_ready         ( DownstreamStackBusLane[34][20].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane20_strm1_cntl          ( DownstreamStackBusLane[34][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane20_strm1_data          ( DownstreamStackBusLane[34][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane20_strm1_data_valid    ( DownstreamStackBusLane[34][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane21_strm0_ready         ( DownstreamStackBusLane[34][21].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane21_strm0_cntl          ( DownstreamStackBusLane[34][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane21_strm0_data          ( DownstreamStackBusLane[34][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane21_strm0_data_valid    ( DownstreamStackBusLane[34][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane21_strm1_ready         ( DownstreamStackBusLane[34][21].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane21_strm1_cntl          ( DownstreamStackBusLane[34][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane21_strm1_data          ( DownstreamStackBusLane[34][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane21_strm1_data_valid    ( DownstreamStackBusLane[34][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane22_strm0_ready         ( DownstreamStackBusLane[34][22].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane22_strm0_cntl          ( DownstreamStackBusLane[34][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane22_strm0_data          ( DownstreamStackBusLane[34][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane22_strm0_data_valid    ( DownstreamStackBusLane[34][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane22_strm1_ready         ( DownstreamStackBusLane[34][22].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane22_strm1_cntl          ( DownstreamStackBusLane[34][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane22_strm1_data          ( DownstreamStackBusLane[34][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane22_strm1_data_valid    ( DownstreamStackBusLane[34][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane23_strm0_ready         ( DownstreamStackBusLane[34][23].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane23_strm0_cntl          ( DownstreamStackBusLane[34][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane23_strm0_data          ( DownstreamStackBusLane[34][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane23_strm0_data_valid    ( DownstreamStackBusLane[34][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane23_strm1_ready         ( DownstreamStackBusLane[34][23].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane23_strm1_cntl          ( DownstreamStackBusLane[34][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane23_strm1_data          ( DownstreamStackBusLane[34][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane23_strm1_data_valid    ( DownstreamStackBusLane[34][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane24_strm0_ready         ( DownstreamStackBusLane[34][24].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane24_strm0_cntl          ( DownstreamStackBusLane[34][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane24_strm0_data          ( DownstreamStackBusLane[34][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane24_strm0_data_valid    ( DownstreamStackBusLane[34][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane24_strm1_ready         ( DownstreamStackBusLane[34][24].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane24_strm1_cntl          ( DownstreamStackBusLane[34][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane24_strm1_data          ( DownstreamStackBusLane[34][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane24_strm1_data_valid    ( DownstreamStackBusLane[34][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane25_strm0_ready         ( DownstreamStackBusLane[34][25].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane25_strm0_cntl          ( DownstreamStackBusLane[34][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane25_strm0_data          ( DownstreamStackBusLane[34][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane25_strm0_data_valid    ( DownstreamStackBusLane[34][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane25_strm1_ready         ( DownstreamStackBusLane[34][25].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane25_strm1_cntl          ( DownstreamStackBusLane[34][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane25_strm1_data          ( DownstreamStackBusLane[34][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane25_strm1_data_valid    ( DownstreamStackBusLane[34][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane26_strm0_ready         ( DownstreamStackBusLane[34][26].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane26_strm0_cntl          ( DownstreamStackBusLane[34][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane26_strm0_data          ( DownstreamStackBusLane[34][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane26_strm0_data_valid    ( DownstreamStackBusLane[34][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane26_strm1_ready         ( DownstreamStackBusLane[34][26].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane26_strm1_cntl          ( DownstreamStackBusLane[34][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane26_strm1_data          ( DownstreamStackBusLane[34][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane26_strm1_data_valid    ( DownstreamStackBusLane[34][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane27_strm0_ready         ( DownstreamStackBusLane[34][27].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane27_strm0_cntl          ( DownstreamStackBusLane[34][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane27_strm0_data          ( DownstreamStackBusLane[34][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane27_strm0_data_valid    ( DownstreamStackBusLane[34][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane27_strm1_ready         ( DownstreamStackBusLane[34][27].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane27_strm1_cntl          ( DownstreamStackBusLane[34][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane27_strm1_data          ( DownstreamStackBusLane[34][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane27_strm1_data_valid    ( DownstreamStackBusLane[34][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane28_strm0_ready         ( DownstreamStackBusLane[34][28].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane28_strm0_cntl          ( DownstreamStackBusLane[34][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane28_strm0_data          ( DownstreamStackBusLane[34][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane28_strm0_data_valid    ( DownstreamStackBusLane[34][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane28_strm1_ready         ( DownstreamStackBusLane[34][28].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane28_strm1_cntl          ( DownstreamStackBusLane[34][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane28_strm1_data          ( DownstreamStackBusLane[34][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane28_strm1_data_valid    ( DownstreamStackBusLane[34][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane29_strm0_ready         ( DownstreamStackBusLane[34][29].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane29_strm0_cntl          ( DownstreamStackBusLane[34][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane29_strm0_data          ( DownstreamStackBusLane[34][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane29_strm0_data_valid    ( DownstreamStackBusLane[34][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane29_strm1_ready         ( DownstreamStackBusLane[34][29].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane29_strm1_cntl          ( DownstreamStackBusLane[34][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane29_strm1_data          ( DownstreamStackBusLane[34][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane29_strm1_data_valid    ( DownstreamStackBusLane[34][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane30_strm0_ready         ( DownstreamStackBusLane[34][30].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane30_strm0_cntl          ( DownstreamStackBusLane[34][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane30_strm0_data          ( DownstreamStackBusLane[34][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane30_strm0_data_valid    ( DownstreamStackBusLane[34][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane30_strm1_ready         ( DownstreamStackBusLane[34][30].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane30_strm1_cntl          ( DownstreamStackBusLane[34][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane30_strm1_data          ( DownstreamStackBusLane[34][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane30_strm1_data_valid    ( DownstreamStackBusLane[34][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 34, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane31_strm0_ready         ( DownstreamStackBusLane[34][31].pe__std__lane_strm0_ready              ),      
        .std__pe34__lane31_strm0_cntl          ( DownstreamStackBusLane[34][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe34__lane31_strm0_data          ( DownstreamStackBusLane[34][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe34__lane31_strm0_data_valid    ( DownstreamStackBusLane[34][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__std__lane31_strm1_ready         ( DownstreamStackBusLane[34][31].pe__std__lane_strm1_ready              ),      
        .std__pe34__lane31_strm1_cntl          ( DownstreamStackBusLane[34][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe34__lane31_strm1_data          ( DownstreamStackBusLane[34][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe34__lane31_strm1_data_valid    ( DownstreamStackBusLane[34][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane0_strm0_ready         ( DownstreamStackBusLane[35][0].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane0_strm0_cntl          ( DownstreamStackBusLane[35][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane0_strm0_data          ( DownstreamStackBusLane[35][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane0_strm0_data_valid    ( DownstreamStackBusLane[35][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane0_strm1_ready         ( DownstreamStackBusLane[35][0].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane0_strm1_cntl          ( DownstreamStackBusLane[35][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane0_strm1_data          ( DownstreamStackBusLane[35][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane0_strm1_data_valid    ( DownstreamStackBusLane[35][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane1_strm0_ready         ( DownstreamStackBusLane[35][1].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane1_strm0_cntl          ( DownstreamStackBusLane[35][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane1_strm0_data          ( DownstreamStackBusLane[35][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane1_strm0_data_valid    ( DownstreamStackBusLane[35][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane1_strm1_ready         ( DownstreamStackBusLane[35][1].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane1_strm1_cntl          ( DownstreamStackBusLane[35][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane1_strm1_data          ( DownstreamStackBusLane[35][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane1_strm1_data_valid    ( DownstreamStackBusLane[35][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane2_strm0_ready         ( DownstreamStackBusLane[35][2].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane2_strm0_cntl          ( DownstreamStackBusLane[35][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane2_strm0_data          ( DownstreamStackBusLane[35][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane2_strm0_data_valid    ( DownstreamStackBusLane[35][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane2_strm1_ready         ( DownstreamStackBusLane[35][2].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane2_strm1_cntl          ( DownstreamStackBusLane[35][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane2_strm1_data          ( DownstreamStackBusLane[35][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane2_strm1_data_valid    ( DownstreamStackBusLane[35][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane3_strm0_ready         ( DownstreamStackBusLane[35][3].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane3_strm0_cntl          ( DownstreamStackBusLane[35][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane3_strm0_data          ( DownstreamStackBusLane[35][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane3_strm0_data_valid    ( DownstreamStackBusLane[35][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane3_strm1_ready         ( DownstreamStackBusLane[35][3].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane3_strm1_cntl          ( DownstreamStackBusLane[35][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane3_strm1_data          ( DownstreamStackBusLane[35][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane3_strm1_data_valid    ( DownstreamStackBusLane[35][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane4_strm0_ready         ( DownstreamStackBusLane[35][4].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane4_strm0_cntl          ( DownstreamStackBusLane[35][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane4_strm0_data          ( DownstreamStackBusLane[35][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane4_strm0_data_valid    ( DownstreamStackBusLane[35][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane4_strm1_ready         ( DownstreamStackBusLane[35][4].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane4_strm1_cntl          ( DownstreamStackBusLane[35][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane4_strm1_data          ( DownstreamStackBusLane[35][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane4_strm1_data_valid    ( DownstreamStackBusLane[35][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane5_strm0_ready         ( DownstreamStackBusLane[35][5].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane5_strm0_cntl          ( DownstreamStackBusLane[35][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane5_strm0_data          ( DownstreamStackBusLane[35][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane5_strm0_data_valid    ( DownstreamStackBusLane[35][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane5_strm1_ready         ( DownstreamStackBusLane[35][5].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane5_strm1_cntl          ( DownstreamStackBusLane[35][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane5_strm1_data          ( DownstreamStackBusLane[35][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane5_strm1_data_valid    ( DownstreamStackBusLane[35][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane6_strm0_ready         ( DownstreamStackBusLane[35][6].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane6_strm0_cntl          ( DownstreamStackBusLane[35][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane6_strm0_data          ( DownstreamStackBusLane[35][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane6_strm0_data_valid    ( DownstreamStackBusLane[35][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane6_strm1_ready         ( DownstreamStackBusLane[35][6].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane6_strm1_cntl          ( DownstreamStackBusLane[35][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane6_strm1_data          ( DownstreamStackBusLane[35][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane6_strm1_data_valid    ( DownstreamStackBusLane[35][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane7_strm0_ready         ( DownstreamStackBusLane[35][7].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane7_strm0_cntl          ( DownstreamStackBusLane[35][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane7_strm0_data          ( DownstreamStackBusLane[35][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane7_strm0_data_valid    ( DownstreamStackBusLane[35][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane7_strm1_ready         ( DownstreamStackBusLane[35][7].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane7_strm1_cntl          ( DownstreamStackBusLane[35][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane7_strm1_data          ( DownstreamStackBusLane[35][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane7_strm1_data_valid    ( DownstreamStackBusLane[35][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane8_strm0_ready         ( DownstreamStackBusLane[35][8].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane8_strm0_cntl          ( DownstreamStackBusLane[35][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane8_strm0_data          ( DownstreamStackBusLane[35][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane8_strm0_data_valid    ( DownstreamStackBusLane[35][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane8_strm1_ready         ( DownstreamStackBusLane[35][8].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane8_strm1_cntl          ( DownstreamStackBusLane[35][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane8_strm1_data          ( DownstreamStackBusLane[35][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane8_strm1_data_valid    ( DownstreamStackBusLane[35][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane9_strm0_ready         ( DownstreamStackBusLane[35][9].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane9_strm0_cntl          ( DownstreamStackBusLane[35][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane9_strm0_data          ( DownstreamStackBusLane[35][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane9_strm0_data_valid    ( DownstreamStackBusLane[35][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane9_strm1_ready         ( DownstreamStackBusLane[35][9].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane9_strm1_cntl          ( DownstreamStackBusLane[35][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane9_strm1_data          ( DownstreamStackBusLane[35][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane9_strm1_data_valid    ( DownstreamStackBusLane[35][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane10_strm0_ready         ( DownstreamStackBusLane[35][10].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane10_strm0_cntl          ( DownstreamStackBusLane[35][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane10_strm0_data          ( DownstreamStackBusLane[35][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane10_strm0_data_valid    ( DownstreamStackBusLane[35][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane10_strm1_ready         ( DownstreamStackBusLane[35][10].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane10_strm1_cntl          ( DownstreamStackBusLane[35][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane10_strm1_data          ( DownstreamStackBusLane[35][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane10_strm1_data_valid    ( DownstreamStackBusLane[35][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane11_strm0_ready         ( DownstreamStackBusLane[35][11].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane11_strm0_cntl          ( DownstreamStackBusLane[35][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane11_strm0_data          ( DownstreamStackBusLane[35][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane11_strm0_data_valid    ( DownstreamStackBusLane[35][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane11_strm1_ready         ( DownstreamStackBusLane[35][11].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane11_strm1_cntl          ( DownstreamStackBusLane[35][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane11_strm1_data          ( DownstreamStackBusLane[35][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane11_strm1_data_valid    ( DownstreamStackBusLane[35][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane12_strm0_ready         ( DownstreamStackBusLane[35][12].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane12_strm0_cntl          ( DownstreamStackBusLane[35][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane12_strm0_data          ( DownstreamStackBusLane[35][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane12_strm0_data_valid    ( DownstreamStackBusLane[35][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane12_strm1_ready         ( DownstreamStackBusLane[35][12].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane12_strm1_cntl          ( DownstreamStackBusLane[35][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane12_strm1_data          ( DownstreamStackBusLane[35][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane12_strm1_data_valid    ( DownstreamStackBusLane[35][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane13_strm0_ready         ( DownstreamStackBusLane[35][13].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane13_strm0_cntl          ( DownstreamStackBusLane[35][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane13_strm0_data          ( DownstreamStackBusLane[35][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane13_strm0_data_valid    ( DownstreamStackBusLane[35][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane13_strm1_ready         ( DownstreamStackBusLane[35][13].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane13_strm1_cntl          ( DownstreamStackBusLane[35][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane13_strm1_data          ( DownstreamStackBusLane[35][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane13_strm1_data_valid    ( DownstreamStackBusLane[35][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane14_strm0_ready         ( DownstreamStackBusLane[35][14].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane14_strm0_cntl          ( DownstreamStackBusLane[35][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane14_strm0_data          ( DownstreamStackBusLane[35][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane14_strm0_data_valid    ( DownstreamStackBusLane[35][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane14_strm1_ready         ( DownstreamStackBusLane[35][14].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane14_strm1_cntl          ( DownstreamStackBusLane[35][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane14_strm1_data          ( DownstreamStackBusLane[35][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane14_strm1_data_valid    ( DownstreamStackBusLane[35][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane15_strm0_ready         ( DownstreamStackBusLane[35][15].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane15_strm0_cntl          ( DownstreamStackBusLane[35][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane15_strm0_data          ( DownstreamStackBusLane[35][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane15_strm0_data_valid    ( DownstreamStackBusLane[35][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane15_strm1_ready         ( DownstreamStackBusLane[35][15].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane15_strm1_cntl          ( DownstreamStackBusLane[35][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane15_strm1_data          ( DownstreamStackBusLane[35][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane15_strm1_data_valid    ( DownstreamStackBusLane[35][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane16_strm0_ready         ( DownstreamStackBusLane[35][16].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane16_strm0_cntl          ( DownstreamStackBusLane[35][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane16_strm0_data          ( DownstreamStackBusLane[35][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane16_strm0_data_valid    ( DownstreamStackBusLane[35][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane16_strm1_ready         ( DownstreamStackBusLane[35][16].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane16_strm1_cntl          ( DownstreamStackBusLane[35][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane16_strm1_data          ( DownstreamStackBusLane[35][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane16_strm1_data_valid    ( DownstreamStackBusLane[35][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane17_strm0_ready         ( DownstreamStackBusLane[35][17].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane17_strm0_cntl          ( DownstreamStackBusLane[35][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane17_strm0_data          ( DownstreamStackBusLane[35][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane17_strm0_data_valid    ( DownstreamStackBusLane[35][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane17_strm1_ready         ( DownstreamStackBusLane[35][17].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane17_strm1_cntl          ( DownstreamStackBusLane[35][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane17_strm1_data          ( DownstreamStackBusLane[35][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane17_strm1_data_valid    ( DownstreamStackBusLane[35][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane18_strm0_ready         ( DownstreamStackBusLane[35][18].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane18_strm0_cntl          ( DownstreamStackBusLane[35][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane18_strm0_data          ( DownstreamStackBusLane[35][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane18_strm0_data_valid    ( DownstreamStackBusLane[35][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane18_strm1_ready         ( DownstreamStackBusLane[35][18].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane18_strm1_cntl          ( DownstreamStackBusLane[35][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane18_strm1_data          ( DownstreamStackBusLane[35][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane18_strm1_data_valid    ( DownstreamStackBusLane[35][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane19_strm0_ready         ( DownstreamStackBusLane[35][19].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane19_strm0_cntl          ( DownstreamStackBusLane[35][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane19_strm0_data          ( DownstreamStackBusLane[35][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane19_strm0_data_valid    ( DownstreamStackBusLane[35][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane19_strm1_ready         ( DownstreamStackBusLane[35][19].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane19_strm1_cntl          ( DownstreamStackBusLane[35][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane19_strm1_data          ( DownstreamStackBusLane[35][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane19_strm1_data_valid    ( DownstreamStackBusLane[35][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane20_strm0_ready         ( DownstreamStackBusLane[35][20].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane20_strm0_cntl          ( DownstreamStackBusLane[35][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane20_strm0_data          ( DownstreamStackBusLane[35][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane20_strm0_data_valid    ( DownstreamStackBusLane[35][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane20_strm1_ready         ( DownstreamStackBusLane[35][20].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane20_strm1_cntl          ( DownstreamStackBusLane[35][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane20_strm1_data          ( DownstreamStackBusLane[35][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane20_strm1_data_valid    ( DownstreamStackBusLane[35][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane21_strm0_ready         ( DownstreamStackBusLane[35][21].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane21_strm0_cntl          ( DownstreamStackBusLane[35][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane21_strm0_data          ( DownstreamStackBusLane[35][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane21_strm0_data_valid    ( DownstreamStackBusLane[35][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane21_strm1_ready         ( DownstreamStackBusLane[35][21].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane21_strm1_cntl          ( DownstreamStackBusLane[35][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane21_strm1_data          ( DownstreamStackBusLane[35][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane21_strm1_data_valid    ( DownstreamStackBusLane[35][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane22_strm0_ready         ( DownstreamStackBusLane[35][22].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane22_strm0_cntl          ( DownstreamStackBusLane[35][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane22_strm0_data          ( DownstreamStackBusLane[35][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane22_strm0_data_valid    ( DownstreamStackBusLane[35][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane22_strm1_ready         ( DownstreamStackBusLane[35][22].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane22_strm1_cntl          ( DownstreamStackBusLane[35][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane22_strm1_data          ( DownstreamStackBusLane[35][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane22_strm1_data_valid    ( DownstreamStackBusLane[35][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane23_strm0_ready         ( DownstreamStackBusLane[35][23].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane23_strm0_cntl          ( DownstreamStackBusLane[35][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane23_strm0_data          ( DownstreamStackBusLane[35][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane23_strm0_data_valid    ( DownstreamStackBusLane[35][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane23_strm1_ready         ( DownstreamStackBusLane[35][23].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane23_strm1_cntl          ( DownstreamStackBusLane[35][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane23_strm1_data          ( DownstreamStackBusLane[35][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane23_strm1_data_valid    ( DownstreamStackBusLane[35][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane24_strm0_ready         ( DownstreamStackBusLane[35][24].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane24_strm0_cntl          ( DownstreamStackBusLane[35][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane24_strm0_data          ( DownstreamStackBusLane[35][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane24_strm0_data_valid    ( DownstreamStackBusLane[35][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane24_strm1_ready         ( DownstreamStackBusLane[35][24].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane24_strm1_cntl          ( DownstreamStackBusLane[35][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane24_strm1_data          ( DownstreamStackBusLane[35][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane24_strm1_data_valid    ( DownstreamStackBusLane[35][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane25_strm0_ready         ( DownstreamStackBusLane[35][25].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane25_strm0_cntl          ( DownstreamStackBusLane[35][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane25_strm0_data          ( DownstreamStackBusLane[35][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane25_strm0_data_valid    ( DownstreamStackBusLane[35][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane25_strm1_ready         ( DownstreamStackBusLane[35][25].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane25_strm1_cntl          ( DownstreamStackBusLane[35][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane25_strm1_data          ( DownstreamStackBusLane[35][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane25_strm1_data_valid    ( DownstreamStackBusLane[35][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane26_strm0_ready         ( DownstreamStackBusLane[35][26].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane26_strm0_cntl          ( DownstreamStackBusLane[35][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane26_strm0_data          ( DownstreamStackBusLane[35][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane26_strm0_data_valid    ( DownstreamStackBusLane[35][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane26_strm1_ready         ( DownstreamStackBusLane[35][26].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane26_strm1_cntl          ( DownstreamStackBusLane[35][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane26_strm1_data          ( DownstreamStackBusLane[35][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane26_strm1_data_valid    ( DownstreamStackBusLane[35][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane27_strm0_ready         ( DownstreamStackBusLane[35][27].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane27_strm0_cntl          ( DownstreamStackBusLane[35][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane27_strm0_data          ( DownstreamStackBusLane[35][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane27_strm0_data_valid    ( DownstreamStackBusLane[35][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane27_strm1_ready         ( DownstreamStackBusLane[35][27].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane27_strm1_cntl          ( DownstreamStackBusLane[35][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane27_strm1_data          ( DownstreamStackBusLane[35][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane27_strm1_data_valid    ( DownstreamStackBusLane[35][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane28_strm0_ready         ( DownstreamStackBusLane[35][28].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane28_strm0_cntl          ( DownstreamStackBusLane[35][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane28_strm0_data          ( DownstreamStackBusLane[35][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane28_strm0_data_valid    ( DownstreamStackBusLane[35][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane28_strm1_ready         ( DownstreamStackBusLane[35][28].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane28_strm1_cntl          ( DownstreamStackBusLane[35][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane28_strm1_data          ( DownstreamStackBusLane[35][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane28_strm1_data_valid    ( DownstreamStackBusLane[35][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane29_strm0_ready         ( DownstreamStackBusLane[35][29].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane29_strm0_cntl          ( DownstreamStackBusLane[35][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane29_strm0_data          ( DownstreamStackBusLane[35][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane29_strm0_data_valid    ( DownstreamStackBusLane[35][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane29_strm1_ready         ( DownstreamStackBusLane[35][29].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane29_strm1_cntl          ( DownstreamStackBusLane[35][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane29_strm1_data          ( DownstreamStackBusLane[35][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane29_strm1_data_valid    ( DownstreamStackBusLane[35][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane30_strm0_ready         ( DownstreamStackBusLane[35][30].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane30_strm0_cntl          ( DownstreamStackBusLane[35][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane30_strm0_data          ( DownstreamStackBusLane[35][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane30_strm0_data_valid    ( DownstreamStackBusLane[35][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane30_strm1_ready         ( DownstreamStackBusLane[35][30].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane30_strm1_cntl          ( DownstreamStackBusLane[35][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane30_strm1_data          ( DownstreamStackBusLane[35][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane30_strm1_data_valid    ( DownstreamStackBusLane[35][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 35, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane31_strm0_ready         ( DownstreamStackBusLane[35][31].pe__std__lane_strm0_ready              ),      
        .std__pe35__lane31_strm0_cntl          ( DownstreamStackBusLane[35][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe35__lane31_strm0_data          ( DownstreamStackBusLane[35][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe35__lane31_strm0_data_valid    ( DownstreamStackBusLane[35][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__std__lane31_strm1_ready         ( DownstreamStackBusLane[35][31].pe__std__lane_strm1_ready              ),      
        .std__pe35__lane31_strm1_cntl          ( DownstreamStackBusLane[35][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe35__lane31_strm1_data          ( DownstreamStackBusLane[35][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe35__lane31_strm1_data_valid    ( DownstreamStackBusLane[35][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane0_strm0_ready         ( DownstreamStackBusLane[36][0].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane0_strm0_cntl          ( DownstreamStackBusLane[36][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane0_strm0_data          ( DownstreamStackBusLane[36][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane0_strm0_data_valid    ( DownstreamStackBusLane[36][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane0_strm1_ready         ( DownstreamStackBusLane[36][0].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane0_strm1_cntl          ( DownstreamStackBusLane[36][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane0_strm1_data          ( DownstreamStackBusLane[36][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane0_strm1_data_valid    ( DownstreamStackBusLane[36][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane1_strm0_ready         ( DownstreamStackBusLane[36][1].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane1_strm0_cntl          ( DownstreamStackBusLane[36][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane1_strm0_data          ( DownstreamStackBusLane[36][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane1_strm0_data_valid    ( DownstreamStackBusLane[36][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane1_strm1_ready         ( DownstreamStackBusLane[36][1].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane1_strm1_cntl          ( DownstreamStackBusLane[36][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane1_strm1_data          ( DownstreamStackBusLane[36][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane1_strm1_data_valid    ( DownstreamStackBusLane[36][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane2_strm0_ready         ( DownstreamStackBusLane[36][2].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane2_strm0_cntl          ( DownstreamStackBusLane[36][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane2_strm0_data          ( DownstreamStackBusLane[36][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane2_strm0_data_valid    ( DownstreamStackBusLane[36][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane2_strm1_ready         ( DownstreamStackBusLane[36][2].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane2_strm1_cntl          ( DownstreamStackBusLane[36][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane2_strm1_data          ( DownstreamStackBusLane[36][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane2_strm1_data_valid    ( DownstreamStackBusLane[36][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane3_strm0_ready         ( DownstreamStackBusLane[36][3].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane3_strm0_cntl          ( DownstreamStackBusLane[36][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane3_strm0_data          ( DownstreamStackBusLane[36][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane3_strm0_data_valid    ( DownstreamStackBusLane[36][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane3_strm1_ready         ( DownstreamStackBusLane[36][3].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane3_strm1_cntl          ( DownstreamStackBusLane[36][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane3_strm1_data          ( DownstreamStackBusLane[36][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane3_strm1_data_valid    ( DownstreamStackBusLane[36][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane4_strm0_ready         ( DownstreamStackBusLane[36][4].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane4_strm0_cntl          ( DownstreamStackBusLane[36][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane4_strm0_data          ( DownstreamStackBusLane[36][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane4_strm0_data_valid    ( DownstreamStackBusLane[36][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane4_strm1_ready         ( DownstreamStackBusLane[36][4].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane4_strm1_cntl          ( DownstreamStackBusLane[36][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane4_strm1_data          ( DownstreamStackBusLane[36][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane4_strm1_data_valid    ( DownstreamStackBusLane[36][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane5_strm0_ready         ( DownstreamStackBusLane[36][5].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane5_strm0_cntl          ( DownstreamStackBusLane[36][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane5_strm0_data          ( DownstreamStackBusLane[36][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane5_strm0_data_valid    ( DownstreamStackBusLane[36][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane5_strm1_ready         ( DownstreamStackBusLane[36][5].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane5_strm1_cntl          ( DownstreamStackBusLane[36][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane5_strm1_data          ( DownstreamStackBusLane[36][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane5_strm1_data_valid    ( DownstreamStackBusLane[36][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane6_strm0_ready         ( DownstreamStackBusLane[36][6].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane6_strm0_cntl          ( DownstreamStackBusLane[36][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane6_strm0_data          ( DownstreamStackBusLane[36][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane6_strm0_data_valid    ( DownstreamStackBusLane[36][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane6_strm1_ready         ( DownstreamStackBusLane[36][6].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane6_strm1_cntl          ( DownstreamStackBusLane[36][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane6_strm1_data          ( DownstreamStackBusLane[36][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane6_strm1_data_valid    ( DownstreamStackBusLane[36][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane7_strm0_ready         ( DownstreamStackBusLane[36][7].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane7_strm0_cntl          ( DownstreamStackBusLane[36][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane7_strm0_data          ( DownstreamStackBusLane[36][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane7_strm0_data_valid    ( DownstreamStackBusLane[36][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane7_strm1_ready         ( DownstreamStackBusLane[36][7].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane7_strm1_cntl          ( DownstreamStackBusLane[36][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane7_strm1_data          ( DownstreamStackBusLane[36][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane7_strm1_data_valid    ( DownstreamStackBusLane[36][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane8_strm0_ready         ( DownstreamStackBusLane[36][8].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane8_strm0_cntl          ( DownstreamStackBusLane[36][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane8_strm0_data          ( DownstreamStackBusLane[36][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane8_strm0_data_valid    ( DownstreamStackBusLane[36][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane8_strm1_ready         ( DownstreamStackBusLane[36][8].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane8_strm1_cntl          ( DownstreamStackBusLane[36][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane8_strm1_data          ( DownstreamStackBusLane[36][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane8_strm1_data_valid    ( DownstreamStackBusLane[36][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane9_strm0_ready         ( DownstreamStackBusLane[36][9].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane9_strm0_cntl          ( DownstreamStackBusLane[36][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane9_strm0_data          ( DownstreamStackBusLane[36][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane9_strm0_data_valid    ( DownstreamStackBusLane[36][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane9_strm1_ready         ( DownstreamStackBusLane[36][9].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane9_strm1_cntl          ( DownstreamStackBusLane[36][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane9_strm1_data          ( DownstreamStackBusLane[36][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane9_strm1_data_valid    ( DownstreamStackBusLane[36][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane10_strm0_ready         ( DownstreamStackBusLane[36][10].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane10_strm0_cntl          ( DownstreamStackBusLane[36][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane10_strm0_data          ( DownstreamStackBusLane[36][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane10_strm0_data_valid    ( DownstreamStackBusLane[36][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane10_strm1_ready         ( DownstreamStackBusLane[36][10].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane10_strm1_cntl          ( DownstreamStackBusLane[36][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane10_strm1_data          ( DownstreamStackBusLane[36][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane10_strm1_data_valid    ( DownstreamStackBusLane[36][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane11_strm0_ready         ( DownstreamStackBusLane[36][11].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane11_strm0_cntl          ( DownstreamStackBusLane[36][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane11_strm0_data          ( DownstreamStackBusLane[36][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane11_strm0_data_valid    ( DownstreamStackBusLane[36][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane11_strm1_ready         ( DownstreamStackBusLane[36][11].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane11_strm1_cntl          ( DownstreamStackBusLane[36][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane11_strm1_data          ( DownstreamStackBusLane[36][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane11_strm1_data_valid    ( DownstreamStackBusLane[36][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane12_strm0_ready         ( DownstreamStackBusLane[36][12].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane12_strm0_cntl          ( DownstreamStackBusLane[36][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane12_strm0_data          ( DownstreamStackBusLane[36][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane12_strm0_data_valid    ( DownstreamStackBusLane[36][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane12_strm1_ready         ( DownstreamStackBusLane[36][12].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane12_strm1_cntl          ( DownstreamStackBusLane[36][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane12_strm1_data          ( DownstreamStackBusLane[36][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane12_strm1_data_valid    ( DownstreamStackBusLane[36][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane13_strm0_ready         ( DownstreamStackBusLane[36][13].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane13_strm0_cntl          ( DownstreamStackBusLane[36][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane13_strm0_data          ( DownstreamStackBusLane[36][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane13_strm0_data_valid    ( DownstreamStackBusLane[36][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane13_strm1_ready         ( DownstreamStackBusLane[36][13].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane13_strm1_cntl          ( DownstreamStackBusLane[36][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane13_strm1_data          ( DownstreamStackBusLane[36][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane13_strm1_data_valid    ( DownstreamStackBusLane[36][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane14_strm0_ready         ( DownstreamStackBusLane[36][14].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane14_strm0_cntl          ( DownstreamStackBusLane[36][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane14_strm0_data          ( DownstreamStackBusLane[36][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane14_strm0_data_valid    ( DownstreamStackBusLane[36][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane14_strm1_ready         ( DownstreamStackBusLane[36][14].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane14_strm1_cntl          ( DownstreamStackBusLane[36][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane14_strm1_data          ( DownstreamStackBusLane[36][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane14_strm1_data_valid    ( DownstreamStackBusLane[36][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane15_strm0_ready         ( DownstreamStackBusLane[36][15].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane15_strm0_cntl          ( DownstreamStackBusLane[36][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane15_strm0_data          ( DownstreamStackBusLane[36][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane15_strm0_data_valid    ( DownstreamStackBusLane[36][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane15_strm1_ready         ( DownstreamStackBusLane[36][15].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane15_strm1_cntl          ( DownstreamStackBusLane[36][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane15_strm1_data          ( DownstreamStackBusLane[36][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane15_strm1_data_valid    ( DownstreamStackBusLane[36][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane16_strm0_ready         ( DownstreamStackBusLane[36][16].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane16_strm0_cntl          ( DownstreamStackBusLane[36][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane16_strm0_data          ( DownstreamStackBusLane[36][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane16_strm0_data_valid    ( DownstreamStackBusLane[36][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane16_strm1_ready         ( DownstreamStackBusLane[36][16].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane16_strm1_cntl          ( DownstreamStackBusLane[36][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane16_strm1_data          ( DownstreamStackBusLane[36][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane16_strm1_data_valid    ( DownstreamStackBusLane[36][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane17_strm0_ready         ( DownstreamStackBusLane[36][17].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane17_strm0_cntl          ( DownstreamStackBusLane[36][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane17_strm0_data          ( DownstreamStackBusLane[36][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane17_strm0_data_valid    ( DownstreamStackBusLane[36][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane17_strm1_ready         ( DownstreamStackBusLane[36][17].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane17_strm1_cntl          ( DownstreamStackBusLane[36][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane17_strm1_data          ( DownstreamStackBusLane[36][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane17_strm1_data_valid    ( DownstreamStackBusLane[36][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane18_strm0_ready         ( DownstreamStackBusLane[36][18].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane18_strm0_cntl          ( DownstreamStackBusLane[36][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane18_strm0_data          ( DownstreamStackBusLane[36][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane18_strm0_data_valid    ( DownstreamStackBusLane[36][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane18_strm1_ready         ( DownstreamStackBusLane[36][18].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane18_strm1_cntl          ( DownstreamStackBusLane[36][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane18_strm1_data          ( DownstreamStackBusLane[36][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane18_strm1_data_valid    ( DownstreamStackBusLane[36][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane19_strm0_ready         ( DownstreamStackBusLane[36][19].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane19_strm0_cntl          ( DownstreamStackBusLane[36][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane19_strm0_data          ( DownstreamStackBusLane[36][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane19_strm0_data_valid    ( DownstreamStackBusLane[36][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane19_strm1_ready         ( DownstreamStackBusLane[36][19].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane19_strm1_cntl          ( DownstreamStackBusLane[36][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane19_strm1_data          ( DownstreamStackBusLane[36][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane19_strm1_data_valid    ( DownstreamStackBusLane[36][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane20_strm0_ready         ( DownstreamStackBusLane[36][20].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane20_strm0_cntl          ( DownstreamStackBusLane[36][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane20_strm0_data          ( DownstreamStackBusLane[36][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane20_strm0_data_valid    ( DownstreamStackBusLane[36][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane20_strm1_ready         ( DownstreamStackBusLane[36][20].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane20_strm1_cntl          ( DownstreamStackBusLane[36][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane20_strm1_data          ( DownstreamStackBusLane[36][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane20_strm1_data_valid    ( DownstreamStackBusLane[36][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane21_strm0_ready         ( DownstreamStackBusLane[36][21].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane21_strm0_cntl          ( DownstreamStackBusLane[36][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane21_strm0_data          ( DownstreamStackBusLane[36][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane21_strm0_data_valid    ( DownstreamStackBusLane[36][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane21_strm1_ready         ( DownstreamStackBusLane[36][21].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane21_strm1_cntl          ( DownstreamStackBusLane[36][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane21_strm1_data          ( DownstreamStackBusLane[36][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane21_strm1_data_valid    ( DownstreamStackBusLane[36][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane22_strm0_ready         ( DownstreamStackBusLane[36][22].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane22_strm0_cntl          ( DownstreamStackBusLane[36][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane22_strm0_data          ( DownstreamStackBusLane[36][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane22_strm0_data_valid    ( DownstreamStackBusLane[36][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane22_strm1_ready         ( DownstreamStackBusLane[36][22].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane22_strm1_cntl          ( DownstreamStackBusLane[36][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane22_strm1_data          ( DownstreamStackBusLane[36][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane22_strm1_data_valid    ( DownstreamStackBusLane[36][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane23_strm0_ready         ( DownstreamStackBusLane[36][23].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane23_strm0_cntl          ( DownstreamStackBusLane[36][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane23_strm0_data          ( DownstreamStackBusLane[36][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane23_strm0_data_valid    ( DownstreamStackBusLane[36][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane23_strm1_ready         ( DownstreamStackBusLane[36][23].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane23_strm1_cntl          ( DownstreamStackBusLane[36][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane23_strm1_data          ( DownstreamStackBusLane[36][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane23_strm1_data_valid    ( DownstreamStackBusLane[36][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane24_strm0_ready         ( DownstreamStackBusLane[36][24].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane24_strm0_cntl          ( DownstreamStackBusLane[36][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane24_strm0_data          ( DownstreamStackBusLane[36][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane24_strm0_data_valid    ( DownstreamStackBusLane[36][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane24_strm1_ready         ( DownstreamStackBusLane[36][24].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane24_strm1_cntl          ( DownstreamStackBusLane[36][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane24_strm1_data          ( DownstreamStackBusLane[36][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane24_strm1_data_valid    ( DownstreamStackBusLane[36][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane25_strm0_ready         ( DownstreamStackBusLane[36][25].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane25_strm0_cntl          ( DownstreamStackBusLane[36][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane25_strm0_data          ( DownstreamStackBusLane[36][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane25_strm0_data_valid    ( DownstreamStackBusLane[36][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane25_strm1_ready         ( DownstreamStackBusLane[36][25].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane25_strm1_cntl          ( DownstreamStackBusLane[36][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane25_strm1_data          ( DownstreamStackBusLane[36][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane25_strm1_data_valid    ( DownstreamStackBusLane[36][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane26_strm0_ready         ( DownstreamStackBusLane[36][26].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane26_strm0_cntl          ( DownstreamStackBusLane[36][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane26_strm0_data          ( DownstreamStackBusLane[36][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane26_strm0_data_valid    ( DownstreamStackBusLane[36][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane26_strm1_ready         ( DownstreamStackBusLane[36][26].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane26_strm1_cntl          ( DownstreamStackBusLane[36][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane26_strm1_data          ( DownstreamStackBusLane[36][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane26_strm1_data_valid    ( DownstreamStackBusLane[36][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane27_strm0_ready         ( DownstreamStackBusLane[36][27].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane27_strm0_cntl          ( DownstreamStackBusLane[36][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane27_strm0_data          ( DownstreamStackBusLane[36][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane27_strm0_data_valid    ( DownstreamStackBusLane[36][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane27_strm1_ready         ( DownstreamStackBusLane[36][27].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane27_strm1_cntl          ( DownstreamStackBusLane[36][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane27_strm1_data          ( DownstreamStackBusLane[36][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane27_strm1_data_valid    ( DownstreamStackBusLane[36][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane28_strm0_ready         ( DownstreamStackBusLane[36][28].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane28_strm0_cntl          ( DownstreamStackBusLane[36][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane28_strm0_data          ( DownstreamStackBusLane[36][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane28_strm0_data_valid    ( DownstreamStackBusLane[36][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane28_strm1_ready         ( DownstreamStackBusLane[36][28].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane28_strm1_cntl          ( DownstreamStackBusLane[36][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane28_strm1_data          ( DownstreamStackBusLane[36][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane28_strm1_data_valid    ( DownstreamStackBusLane[36][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane29_strm0_ready         ( DownstreamStackBusLane[36][29].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane29_strm0_cntl          ( DownstreamStackBusLane[36][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane29_strm0_data          ( DownstreamStackBusLane[36][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane29_strm0_data_valid    ( DownstreamStackBusLane[36][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane29_strm1_ready         ( DownstreamStackBusLane[36][29].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane29_strm1_cntl          ( DownstreamStackBusLane[36][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane29_strm1_data          ( DownstreamStackBusLane[36][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane29_strm1_data_valid    ( DownstreamStackBusLane[36][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane30_strm0_ready         ( DownstreamStackBusLane[36][30].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane30_strm0_cntl          ( DownstreamStackBusLane[36][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane30_strm0_data          ( DownstreamStackBusLane[36][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane30_strm0_data_valid    ( DownstreamStackBusLane[36][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane30_strm1_ready         ( DownstreamStackBusLane[36][30].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane30_strm1_cntl          ( DownstreamStackBusLane[36][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane30_strm1_data          ( DownstreamStackBusLane[36][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane30_strm1_data_valid    ( DownstreamStackBusLane[36][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 36, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane31_strm0_ready         ( DownstreamStackBusLane[36][31].pe__std__lane_strm0_ready              ),      
        .std__pe36__lane31_strm0_cntl          ( DownstreamStackBusLane[36][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe36__lane31_strm0_data          ( DownstreamStackBusLane[36][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe36__lane31_strm0_data_valid    ( DownstreamStackBusLane[36][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__std__lane31_strm1_ready         ( DownstreamStackBusLane[36][31].pe__std__lane_strm1_ready              ),      
        .std__pe36__lane31_strm1_cntl          ( DownstreamStackBusLane[36][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe36__lane31_strm1_data          ( DownstreamStackBusLane[36][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe36__lane31_strm1_data_valid    ( DownstreamStackBusLane[36][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane0_strm0_ready         ( DownstreamStackBusLane[37][0].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane0_strm0_cntl          ( DownstreamStackBusLane[37][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane0_strm0_data          ( DownstreamStackBusLane[37][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane0_strm0_data_valid    ( DownstreamStackBusLane[37][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane0_strm1_ready         ( DownstreamStackBusLane[37][0].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane0_strm1_cntl          ( DownstreamStackBusLane[37][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane0_strm1_data          ( DownstreamStackBusLane[37][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane0_strm1_data_valid    ( DownstreamStackBusLane[37][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane1_strm0_ready         ( DownstreamStackBusLane[37][1].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane1_strm0_cntl          ( DownstreamStackBusLane[37][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane1_strm0_data          ( DownstreamStackBusLane[37][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane1_strm0_data_valid    ( DownstreamStackBusLane[37][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane1_strm1_ready         ( DownstreamStackBusLane[37][1].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane1_strm1_cntl          ( DownstreamStackBusLane[37][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane1_strm1_data          ( DownstreamStackBusLane[37][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane1_strm1_data_valid    ( DownstreamStackBusLane[37][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane2_strm0_ready         ( DownstreamStackBusLane[37][2].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane2_strm0_cntl          ( DownstreamStackBusLane[37][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane2_strm0_data          ( DownstreamStackBusLane[37][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane2_strm0_data_valid    ( DownstreamStackBusLane[37][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane2_strm1_ready         ( DownstreamStackBusLane[37][2].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane2_strm1_cntl          ( DownstreamStackBusLane[37][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane2_strm1_data          ( DownstreamStackBusLane[37][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane2_strm1_data_valid    ( DownstreamStackBusLane[37][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane3_strm0_ready         ( DownstreamStackBusLane[37][3].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane3_strm0_cntl          ( DownstreamStackBusLane[37][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane3_strm0_data          ( DownstreamStackBusLane[37][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane3_strm0_data_valid    ( DownstreamStackBusLane[37][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane3_strm1_ready         ( DownstreamStackBusLane[37][3].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane3_strm1_cntl          ( DownstreamStackBusLane[37][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane3_strm1_data          ( DownstreamStackBusLane[37][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane3_strm1_data_valid    ( DownstreamStackBusLane[37][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane4_strm0_ready         ( DownstreamStackBusLane[37][4].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane4_strm0_cntl          ( DownstreamStackBusLane[37][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane4_strm0_data          ( DownstreamStackBusLane[37][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane4_strm0_data_valid    ( DownstreamStackBusLane[37][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane4_strm1_ready         ( DownstreamStackBusLane[37][4].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane4_strm1_cntl          ( DownstreamStackBusLane[37][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane4_strm1_data          ( DownstreamStackBusLane[37][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane4_strm1_data_valid    ( DownstreamStackBusLane[37][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane5_strm0_ready         ( DownstreamStackBusLane[37][5].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane5_strm0_cntl          ( DownstreamStackBusLane[37][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane5_strm0_data          ( DownstreamStackBusLane[37][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane5_strm0_data_valid    ( DownstreamStackBusLane[37][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane5_strm1_ready         ( DownstreamStackBusLane[37][5].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane5_strm1_cntl          ( DownstreamStackBusLane[37][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane5_strm1_data          ( DownstreamStackBusLane[37][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane5_strm1_data_valid    ( DownstreamStackBusLane[37][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane6_strm0_ready         ( DownstreamStackBusLane[37][6].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane6_strm0_cntl          ( DownstreamStackBusLane[37][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane6_strm0_data          ( DownstreamStackBusLane[37][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane6_strm0_data_valid    ( DownstreamStackBusLane[37][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane6_strm1_ready         ( DownstreamStackBusLane[37][6].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane6_strm1_cntl          ( DownstreamStackBusLane[37][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane6_strm1_data          ( DownstreamStackBusLane[37][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane6_strm1_data_valid    ( DownstreamStackBusLane[37][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane7_strm0_ready         ( DownstreamStackBusLane[37][7].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane7_strm0_cntl          ( DownstreamStackBusLane[37][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane7_strm0_data          ( DownstreamStackBusLane[37][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane7_strm0_data_valid    ( DownstreamStackBusLane[37][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane7_strm1_ready         ( DownstreamStackBusLane[37][7].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane7_strm1_cntl          ( DownstreamStackBusLane[37][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane7_strm1_data          ( DownstreamStackBusLane[37][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane7_strm1_data_valid    ( DownstreamStackBusLane[37][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane8_strm0_ready         ( DownstreamStackBusLane[37][8].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane8_strm0_cntl          ( DownstreamStackBusLane[37][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane8_strm0_data          ( DownstreamStackBusLane[37][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane8_strm0_data_valid    ( DownstreamStackBusLane[37][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane8_strm1_ready         ( DownstreamStackBusLane[37][8].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane8_strm1_cntl          ( DownstreamStackBusLane[37][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane8_strm1_data          ( DownstreamStackBusLane[37][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane8_strm1_data_valid    ( DownstreamStackBusLane[37][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane9_strm0_ready         ( DownstreamStackBusLane[37][9].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane9_strm0_cntl          ( DownstreamStackBusLane[37][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane9_strm0_data          ( DownstreamStackBusLane[37][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane9_strm0_data_valid    ( DownstreamStackBusLane[37][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane9_strm1_ready         ( DownstreamStackBusLane[37][9].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane9_strm1_cntl          ( DownstreamStackBusLane[37][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane9_strm1_data          ( DownstreamStackBusLane[37][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane9_strm1_data_valid    ( DownstreamStackBusLane[37][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane10_strm0_ready         ( DownstreamStackBusLane[37][10].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane10_strm0_cntl          ( DownstreamStackBusLane[37][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane10_strm0_data          ( DownstreamStackBusLane[37][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane10_strm0_data_valid    ( DownstreamStackBusLane[37][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane10_strm1_ready         ( DownstreamStackBusLane[37][10].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane10_strm1_cntl          ( DownstreamStackBusLane[37][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane10_strm1_data          ( DownstreamStackBusLane[37][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane10_strm1_data_valid    ( DownstreamStackBusLane[37][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane11_strm0_ready         ( DownstreamStackBusLane[37][11].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane11_strm0_cntl          ( DownstreamStackBusLane[37][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane11_strm0_data          ( DownstreamStackBusLane[37][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane11_strm0_data_valid    ( DownstreamStackBusLane[37][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane11_strm1_ready         ( DownstreamStackBusLane[37][11].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane11_strm1_cntl          ( DownstreamStackBusLane[37][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane11_strm1_data          ( DownstreamStackBusLane[37][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane11_strm1_data_valid    ( DownstreamStackBusLane[37][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane12_strm0_ready         ( DownstreamStackBusLane[37][12].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane12_strm0_cntl          ( DownstreamStackBusLane[37][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane12_strm0_data          ( DownstreamStackBusLane[37][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane12_strm0_data_valid    ( DownstreamStackBusLane[37][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane12_strm1_ready         ( DownstreamStackBusLane[37][12].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane12_strm1_cntl          ( DownstreamStackBusLane[37][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane12_strm1_data          ( DownstreamStackBusLane[37][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane12_strm1_data_valid    ( DownstreamStackBusLane[37][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane13_strm0_ready         ( DownstreamStackBusLane[37][13].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane13_strm0_cntl          ( DownstreamStackBusLane[37][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane13_strm0_data          ( DownstreamStackBusLane[37][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane13_strm0_data_valid    ( DownstreamStackBusLane[37][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane13_strm1_ready         ( DownstreamStackBusLane[37][13].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane13_strm1_cntl          ( DownstreamStackBusLane[37][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane13_strm1_data          ( DownstreamStackBusLane[37][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane13_strm1_data_valid    ( DownstreamStackBusLane[37][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane14_strm0_ready         ( DownstreamStackBusLane[37][14].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane14_strm0_cntl          ( DownstreamStackBusLane[37][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane14_strm0_data          ( DownstreamStackBusLane[37][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane14_strm0_data_valid    ( DownstreamStackBusLane[37][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane14_strm1_ready         ( DownstreamStackBusLane[37][14].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane14_strm1_cntl          ( DownstreamStackBusLane[37][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane14_strm1_data          ( DownstreamStackBusLane[37][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane14_strm1_data_valid    ( DownstreamStackBusLane[37][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane15_strm0_ready         ( DownstreamStackBusLane[37][15].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane15_strm0_cntl          ( DownstreamStackBusLane[37][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane15_strm0_data          ( DownstreamStackBusLane[37][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane15_strm0_data_valid    ( DownstreamStackBusLane[37][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane15_strm1_ready         ( DownstreamStackBusLane[37][15].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane15_strm1_cntl          ( DownstreamStackBusLane[37][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane15_strm1_data          ( DownstreamStackBusLane[37][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane15_strm1_data_valid    ( DownstreamStackBusLane[37][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane16_strm0_ready         ( DownstreamStackBusLane[37][16].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane16_strm0_cntl          ( DownstreamStackBusLane[37][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane16_strm0_data          ( DownstreamStackBusLane[37][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane16_strm0_data_valid    ( DownstreamStackBusLane[37][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane16_strm1_ready         ( DownstreamStackBusLane[37][16].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane16_strm1_cntl          ( DownstreamStackBusLane[37][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane16_strm1_data          ( DownstreamStackBusLane[37][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane16_strm1_data_valid    ( DownstreamStackBusLane[37][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane17_strm0_ready         ( DownstreamStackBusLane[37][17].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane17_strm0_cntl          ( DownstreamStackBusLane[37][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane17_strm0_data          ( DownstreamStackBusLane[37][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane17_strm0_data_valid    ( DownstreamStackBusLane[37][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane17_strm1_ready         ( DownstreamStackBusLane[37][17].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane17_strm1_cntl          ( DownstreamStackBusLane[37][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane17_strm1_data          ( DownstreamStackBusLane[37][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane17_strm1_data_valid    ( DownstreamStackBusLane[37][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane18_strm0_ready         ( DownstreamStackBusLane[37][18].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane18_strm0_cntl          ( DownstreamStackBusLane[37][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane18_strm0_data          ( DownstreamStackBusLane[37][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane18_strm0_data_valid    ( DownstreamStackBusLane[37][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane18_strm1_ready         ( DownstreamStackBusLane[37][18].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane18_strm1_cntl          ( DownstreamStackBusLane[37][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane18_strm1_data          ( DownstreamStackBusLane[37][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane18_strm1_data_valid    ( DownstreamStackBusLane[37][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane19_strm0_ready         ( DownstreamStackBusLane[37][19].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane19_strm0_cntl          ( DownstreamStackBusLane[37][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane19_strm0_data          ( DownstreamStackBusLane[37][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane19_strm0_data_valid    ( DownstreamStackBusLane[37][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane19_strm1_ready         ( DownstreamStackBusLane[37][19].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane19_strm1_cntl          ( DownstreamStackBusLane[37][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane19_strm1_data          ( DownstreamStackBusLane[37][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane19_strm1_data_valid    ( DownstreamStackBusLane[37][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane20_strm0_ready         ( DownstreamStackBusLane[37][20].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane20_strm0_cntl          ( DownstreamStackBusLane[37][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane20_strm0_data          ( DownstreamStackBusLane[37][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane20_strm0_data_valid    ( DownstreamStackBusLane[37][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane20_strm1_ready         ( DownstreamStackBusLane[37][20].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane20_strm1_cntl          ( DownstreamStackBusLane[37][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane20_strm1_data          ( DownstreamStackBusLane[37][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane20_strm1_data_valid    ( DownstreamStackBusLane[37][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane21_strm0_ready         ( DownstreamStackBusLane[37][21].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane21_strm0_cntl          ( DownstreamStackBusLane[37][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane21_strm0_data          ( DownstreamStackBusLane[37][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane21_strm0_data_valid    ( DownstreamStackBusLane[37][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane21_strm1_ready         ( DownstreamStackBusLane[37][21].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane21_strm1_cntl          ( DownstreamStackBusLane[37][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane21_strm1_data          ( DownstreamStackBusLane[37][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane21_strm1_data_valid    ( DownstreamStackBusLane[37][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane22_strm0_ready         ( DownstreamStackBusLane[37][22].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane22_strm0_cntl          ( DownstreamStackBusLane[37][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane22_strm0_data          ( DownstreamStackBusLane[37][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane22_strm0_data_valid    ( DownstreamStackBusLane[37][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane22_strm1_ready         ( DownstreamStackBusLane[37][22].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane22_strm1_cntl          ( DownstreamStackBusLane[37][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane22_strm1_data          ( DownstreamStackBusLane[37][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane22_strm1_data_valid    ( DownstreamStackBusLane[37][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane23_strm0_ready         ( DownstreamStackBusLane[37][23].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane23_strm0_cntl          ( DownstreamStackBusLane[37][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane23_strm0_data          ( DownstreamStackBusLane[37][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane23_strm0_data_valid    ( DownstreamStackBusLane[37][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane23_strm1_ready         ( DownstreamStackBusLane[37][23].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane23_strm1_cntl          ( DownstreamStackBusLane[37][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane23_strm1_data          ( DownstreamStackBusLane[37][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane23_strm1_data_valid    ( DownstreamStackBusLane[37][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane24_strm0_ready         ( DownstreamStackBusLane[37][24].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane24_strm0_cntl          ( DownstreamStackBusLane[37][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane24_strm0_data          ( DownstreamStackBusLane[37][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane24_strm0_data_valid    ( DownstreamStackBusLane[37][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane24_strm1_ready         ( DownstreamStackBusLane[37][24].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane24_strm1_cntl          ( DownstreamStackBusLane[37][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane24_strm1_data          ( DownstreamStackBusLane[37][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane24_strm1_data_valid    ( DownstreamStackBusLane[37][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane25_strm0_ready         ( DownstreamStackBusLane[37][25].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane25_strm0_cntl          ( DownstreamStackBusLane[37][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane25_strm0_data          ( DownstreamStackBusLane[37][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane25_strm0_data_valid    ( DownstreamStackBusLane[37][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane25_strm1_ready         ( DownstreamStackBusLane[37][25].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane25_strm1_cntl          ( DownstreamStackBusLane[37][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane25_strm1_data          ( DownstreamStackBusLane[37][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane25_strm1_data_valid    ( DownstreamStackBusLane[37][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane26_strm0_ready         ( DownstreamStackBusLane[37][26].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane26_strm0_cntl          ( DownstreamStackBusLane[37][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane26_strm0_data          ( DownstreamStackBusLane[37][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane26_strm0_data_valid    ( DownstreamStackBusLane[37][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane26_strm1_ready         ( DownstreamStackBusLane[37][26].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane26_strm1_cntl          ( DownstreamStackBusLane[37][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane26_strm1_data          ( DownstreamStackBusLane[37][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane26_strm1_data_valid    ( DownstreamStackBusLane[37][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane27_strm0_ready         ( DownstreamStackBusLane[37][27].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane27_strm0_cntl          ( DownstreamStackBusLane[37][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane27_strm0_data          ( DownstreamStackBusLane[37][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane27_strm0_data_valid    ( DownstreamStackBusLane[37][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane27_strm1_ready         ( DownstreamStackBusLane[37][27].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane27_strm1_cntl          ( DownstreamStackBusLane[37][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane27_strm1_data          ( DownstreamStackBusLane[37][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane27_strm1_data_valid    ( DownstreamStackBusLane[37][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane28_strm0_ready         ( DownstreamStackBusLane[37][28].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane28_strm0_cntl          ( DownstreamStackBusLane[37][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane28_strm0_data          ( DownstreamStackBusLane[37][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane28_strm0_data_valid    ( DownstreamStackBusLane[37][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane28_strm1_ready         ( DownstreamStackBusLane[37][28].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane28_strm1_cntl          ( DownstreamStackBusLane[37][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane28_strm1_data          ( DownstreamStackBusLane[37][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane28_strm1_data_valid    ( DownstreamStackBusLane[37][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane29_strm0_ready         ( DownstreamStackBusLane[37][29].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane29_strm0_cntl          ( DownstreamStackBusLane[37][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane29_strm0_data          ( DownstreamStackBusLane[37][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane29_strm0_data_valid    ( DownstreamStackBusLane[37][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane29_strm1_ready         ( DownstreamStackBusLane[37][29].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane29_strm1_cntl          ( DownstreamStackBusLane[37][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane29_strm1_data          ( DownstreamStackBusLane[37][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane29_strm1_data_valid    ( DownstreamStackBusLane[37][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane30_strm0_ready         ( DownstreamStackBusLane[37][30].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane30_strm0_cntl          ( DownstreamStackBusLane[37][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane30_strm0_data          ( DownstreamStackBusLane[37][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane30_strm0_data_valid    ( DownstreamStackBusLane[37][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane30_strm1_ready         ( DownstreamStackBusLane[37][30].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane30_strm1_cntl          ( DownstreamStackBusLane[37][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane30_strm1_data          ( DownstreamStackBusLane[37][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane30_strm1_data_valid    ( DownstreamStackBusLane[37][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 37, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane31_strm0_ready         ( DownstreamStackBusLane[37][31].pe__std__lane_strm0_ready              ),      
        .std__pe37__lane31_strm0_cntl          ( DownstreamStackBusLane[37][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe37__lane31_strm0_data          ( DownstreamStackBusLane[37][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe37__lane31_strm0_data_valid    ( DownstreamStackBusLane[37][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__std__lane31_strm1_ready         ( DownstreamStackBusLane[37][31].pe__std__lane_strm1_ready              ),      
        .std__pe37__lane31_strm1_cntl          ( DownstreamStackBusLane[37][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe37__lane31_strm1_data          ( DownstreamStackBusLane[37][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe37__lane31_strm1_data_valid    ( DownstreamStackBusLane[37][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane0_strm0_ready         ( DownstreamStackBusLane[38][0].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane0_strm0_cntl          ( DownstreamStackBusLane[38][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane0_strm0_data          ( DownstreamStackBusLane[38][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane0_strm0_data_valid    ( DownstreamStackBusLane[38][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane0_strm1_ready         ( DownstreamStackBusLane[38][0].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane0_strm1_cntl          ( DownstreamStackBusLane[38][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane0_strm1_data          ( DownstreamStackBusLane[38][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane0_strm1_data_valid    ( DownstreamStackBusLane[38][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane1_strm0_ready         ( DownstreamStackBusLane[38][1].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane1_strm0_cntl          ( DownstreamStackBusLane[38][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane1_strm0_data          ( DownstreamStackBusLane[38][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane1_strm0_data_valid    ( DownstreamStackBusLane[38][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane1_strm1_ready         ( DownstreamStackBusLane[38][1].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane1_strm1_cntl          ( DownstreamStackBusLane[38][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane1_strm1_data          ( DownstreamStackBusLane[38][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane1_strm1_data_valid    ( DownstreamStackBusLane[38][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane2_strm0_ready         ( DownstreamStackBusLane[38][2].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane2_strm0_cntl          ( DownstreamStackBusLane[38][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane2_strm0_data          ( DownstreamStackBusLane[38][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane2_strm0_data_valid    ( DownstreamStackBusLane[38][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane2_strm1_ready         ( DownstreamStackBusLane[38][2].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane2_strm1_cntl          ( DownstreamStackBusLane[38][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane2_strm1_data          ( DownstreamStackBusLane[38][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane2_strm1_data_valid    ( DownstreamStackBusLane[38][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane3_strm0_ready         ( DownstreamStackBusLane[38][3].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane3_strm0_cntl          ( DownstreamStackBusLane[38][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane3_strm0_data          ( DownstreamStackBusLane[38][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane3_strm0_data_valid    ( DownstreamStackBusLane[38][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane3_strm1_ready         ( DownstreamStackBusLane[38][3].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane3_strm1_cntl          ( DownstreamStackBusLane[38][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane3_strm1_data          ( DownstreamStackBusLane[38][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane3_strm1_data_valid    ( DownstreamStackBusLane[38][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane4_strm0_ready         ( DownstreamStackBusLane[38][4].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane4_strm0_cntl          ( DownstreamStackBusLane[38][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane4_strm0_data          ( DownstreamStackBusLane[38][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane4_strm0_data_valid    ( DownstreamStackBusLane[38][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane4_strm1_ready         ( DownstreamStackBusLane[38][4].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane4_strm1_cntl          ( DownstreamStackBusLane[38][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane4_strm1_data          ( DownstreamStackBusLane[38][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane4_strm1_data_valid    ( DownstreamStackBusLane[38][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane5_strm0_ready         ( DownstreamStackBusLane[38][5].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane5_strm0_cntl          ( DownstreamStackBusLane[38][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane5_strm0_data          ( DownstreamStackBusLane[38][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane5_strm0_data_valid    ( DownstreamStackBusLane[38][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane5_strm1_ready         ( DownstreamStackBusLane[38][5].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane5_strm1_cntl          ( DownstreamStackBusLane[38][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane5_strm1_data          ( DownstreamStackBusLane[38][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane5_strm1_data_valid    ( DownstreamStackBusLane[38][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane6_strm0_ready         ( DownstreamStackBusLane[38][6].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane6_strm0_cntl          ( DownstreamStackBusLane[38][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane6_strm0_data          ( DownstreamStackBusLane[38][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane6_strm0_data_valid    ( DownstreamStackBusLane[38][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane6_strm1_ready         ( DownstreamStackBusLane[38][6].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane6_strm1_cntl          ( DownstreamStackBusLane[38][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane6_strm1_data          ( DownstreamStackBusLane[38][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane6_strm1_data_valid    ( DownstreamStackBusLane[38][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane7_strm0_ready         ( DownstreamStackBusLane[38][7].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane7_strm0_cntl          ( DownstreamStackBusLane[38][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane7_strm0_data          ( DownstreamStackBusLane[38][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane7_strm0_data_valid    ( DownstreamStackBusLane[38][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane7_strm1_ready         ( DownstreamStackBusLane[38][7].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane7_strm1_cntl          ( DownstreamStackBusLane[38][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane7_strm1_data          ( DownstreamStackBusLane[38][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane7_strm1_data_valid    ( DownstreamStackBusLane[38][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane8_strm0_ready         ( DownstreamStackBusLane[38][8].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane8_strm0_cntl          ( DownstreamStackBusLane[38][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane8_strm0_data          ( DownstreamStackBusLane[38][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane8_strm0_data_valid    ( DownstreamStackBusLane[38][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane8_strm1_ready         ( DownstreamStackBusLane[38][8].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane8_strm1_cntl          ( DownstreamStackBusLane[38][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane8_strm1_data          ( DownstreamStackBusLane[38][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane8_strm1_data_valid    ( DownstreamStackBusLane[38][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane9_strm0_ready         ( DownstreamStackBusLane[38][9].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane9_strm0_cntl          ( DownstreamStackBusLane[38][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane9_strm0_data          ( DownstreamStackBusLane[38][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane9_strm0_data_valid    ( DownstreamStackBusLane[38][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane9_strm1_ready         ( DownstreamStackBusLane[38][9].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane9_strm1_cntl          ( DownstreamStackBusLane[38][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane9_strm1_data          ( DownstreamStackBusLane[38][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane9_strm1_data_valid    ( DownstreamStackBusLane[38][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane10_strm0_ready         ( DownstreamStackBusLane[38][10].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane10_strm0_cntl          ( DownstreamStackBusLane[38][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane10_strm0_data          ( DownstreamStackBusLane[38][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane10_strm0_data_valid    ( DownstreamStackBusLane[38][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane10_strm1_ready         ( DownstreamStackBusLane[38][10].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane10_strm1_cntl          ( DownstreamStackBusLane[38][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane10_strm1_data          ( DownstreamStackBusLane[38][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane10_strm1_data_valid    ( DownstreamStackBusLane[38][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane11_strm0_ready         ( DownstreamStackBusLane[38][11].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane11_strm0_cntl          ( DownstreamStackBusLane[38][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane11_strm0_data          ( DownstreamStackBusLane[38][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane11_strm0_data_valid    ( DownstreamStackBusLane[38][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane11_strm1_ready         ( DownstreamStackBusLane[38][11].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane11_strm1_cntl          ( DownstreamStackBusLane[38][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane11_strm1_data          ( DownstreamStackBusLane[38][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane11_strm1_data_valid    ( DownstreamStackBusLane[38][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane12_strm0_ready         ( DownstreamStackBusLane[38][12].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane12_strm0_cntl          ( DownstreamStackBusLane[38][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane12_strm0_data          ( DownstreamStackBusLane[38][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane12_strm0_data_valid    ( DownstreamStackBusLane[38][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane12_strm1_ready         ( DownstreamStackBusLane[38][12].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane12_strm1_cntl          ( DownstreamStackBusLane[38][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane12_strm1_data          ( DownstreamStackBusLane[38][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane12_strm1_data_valid    ( DownstreamStackBusLane[38][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane13_strm0_ready         ( DownstreamStackBusLane[38][13].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane13_strm0_cntl          ( DownstreamStackBusLane[38][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane13_strm0_data          ( DownstreamStackBusLane[38][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane13_strm0_data_valid    ( DownstreamStackBusLane[38][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane13_strm1_ready         ( DownstreamStackBusLane[38][13].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane13_strm1_cntl          ( DownstreamStackBusLane[38][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane13_strm1_data          ( DownstreamStackBusLane[38][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane13_strm1_data_valid    ( DownstreamStackBusLane[38][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane14_strm0_ready         ( DownstreamStackBusLane[38][14].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane14_strm0_cntl          ( DownstreamStackBusLane[38][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane14_strm0_data          ( DownstreamStackBusLane[38][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane14_strm0_data_valid    ( DownstreamStackBusLane[38][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane14_strm1_ready         ( DownstreamStackBusLane[38][14].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane14_strm1_cntl          ( DownstreamStackBusLane[38][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane14_strm1_data          ( DownstreamStackBusLane[38][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane14_strm1_data_valid    ( DownstreamStackBusLane[38][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane15_strm0_ready         ( DownstreamStackBusLane[38][15].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane15_strm0_cntl          ( DownstreamStackBusLane[38][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane15_strm0_data          ( DownstreamStackBusLane[38][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane15_strm0_data_valid    ( DownstreamStackBusLane[38][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane15_strm1_ready         ( DownstreamStackBusLane[38][15].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane15_strm1_cntl          ( DownstreamStackBusLane[38][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane15_strm1_data          ( DownstreamStackBusLane[38][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane15_strm1_data_valid    ( DownstreamStackBusLane[38][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane16_strm0_ready         ( DownstreamStackBusLane[38][16].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane16_strm0_cntl          ( DownstreamStackBusLane[38][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane16_strm0_data          ( DownstreamStackBusLane[38][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane16_strm0_data_valid    ( DownstreamStackBusLane[38][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane16_strm1_ready         ( DownstreamStackBusLane[38][16].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane16_strm1_cntl          ( DownstreamStackBusLane[38][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane16_strm1_data          ( DownstreamStackBusLane[38][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane16_strm1_data_valid    ( DownstreamStackBusLane[38][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane17_strm0_ready         ( DownstreamStackBusLane[38][17].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane17_strm0_cntl          ( DownstreamStackBusLane[38][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane17_strm0_data          ( DownstreamStackBusLane[38][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane17_strm0_data_valid    ( DownstreamStackBusLane[38][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane17_strm1_ready         ( DownstreamStackBusLane[38][17].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane17_strm1_cntl          ( DownstreamStackBusLane[38][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane17_strm1_data          ( DownstreamStackBusLane[38][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane17_strm1_data_valid    ( DownstreamStackBusLane[38][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane18_strm0_ready         ( DownstreamStackBusLane[38][18].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane18_strm0_cntl          ( DownstreamStackBusLane[38][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane18_strm0_data          ( DownstreamStackBusLane[38][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane18_strm0_data_valid    ( DownstreamStackBusLane[38][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane18_strm1_ready         ( DownstreamStackBusLane[38][18].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane18_strm1_cntl          ( DownstreamStackBusLane[38][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane18_strm1_data          ( DownstreamStackBusLane[38][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane18_strm1_data_valid    ( DownstreamStackBusLane[38][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane19_strm0_ready         ( DownstreamStackBusLane[38][19].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane19_strm0_cntl          ( DownstreamStackBusLane[38][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane19_strm0_data          ( DownstreamStackBusLane[38][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane19_strm0_data_valid    ( DownstreamStackBusLane[38][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane19_strm1_ready         ( DownstreamStackBusLane[38][19].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane19_strm1_cntl          ( DownstreamStackBusLane[38][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane19_strm1_data          ( DownstreamStackBusLane[38][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane19_strm1_data_valid    ( DownstreamStackBusLane[38][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane20_strm0_ready         ( DownstreamStackBusLane[38][20].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane20_strm0_cntl          ( DownstreamStackBusLane[38][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane20_strm0_data          ( DownstreamStackBusLane[38][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane20_strm0_data_valid    ( DownstreamStackBusLane[38][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane20_strm1_ready         ( DownstreamStackBusLane[38][20].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane20_strm1_cntl          ( DownstreamStackBusLane[38][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane20_strm1_data          ( DownstreamStackBusLane[38][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane20_strm1_data_valid    ( DownstreamStackBusLane[38][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane21_strm0_ready         ( DownstreamStackBusLane[38][21].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane21_strm0_cntl          ( DownstreamStackBusLane[38][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane21_strm0_data          ( DownstreamStackBusLane[38][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane21_strm0_data_valid    ( DownstreamStackBusLane[38][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane21_strm1_ready         ( DownstreamStackBusLane[38][21].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane21_strm1_cntl          ( DownstreamStackBusLane[38][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane21_strm1_data          ( DownstreamStackBusLane[38][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane21_strm1_data_valid    ( DownstreamStackBusLane[38][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane22_strm0_ready         ( DownstreamStackBusLane[38][22].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane22_strm0_cntl          ( DownstreamStackBusLane[38][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane22_strm0_data          ( DownstreamStackBusLane[38][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane22_strm0_data_valid    ( DownstreamStackBusLane[38][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane22_strm1_ready         ( DownstreamStackBusLane[38][22].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane22_strm1_cntl          ( DownstreamStackBusLane[38][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane22_strm1_data          ( DownstreamStackBusLane[38][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane22_strm1_data_valid    ( DownstreamStackBusLane[38][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane23_strm0_ready         ( DownstreamStackBusLane[38][23].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane23_strm0_cntl          ( DownstreamStackBusLane[38][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane23_strm0_data          ( DownstreamStackBusLane[38][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane23_strm0_data_valid    ( DownstreamStackBusLane[38][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane23_strm1_ready         ( DownstreamStackBusLane[38][23].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane23_strm1_cntl          ( DownstreamStackBusLane[38][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane23_strm1_data          ( DownstreamStackBusLane[38][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane23_strm1_data_valid    ( DownstreamStackBusLane[38][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane24_strm0_ready         ( DownstreamStackBusLane[38][24].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane24_strm0_cntl          ( DownstreamStackBusLane[38][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane24_strm0_data          ( DownstreamStackBusLane[38][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane24_strm0_data_valid    ( DownstreamStackBusLane[38][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane24_strm1_ready         ( DownstreamStackBusLane[38][24].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane24_strm1_cntl          ( DownstreamStackBusLane[38][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane24_strm1_data          ( DownstreamStackBusLane[38][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane24_strm1_data_valid    ( DownstreamStackBusLane[38][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane25_strm0_ready         ( DownstreamStackBusLane[38][25].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane25_strm0_cntl          ( DownstreamStackBusLane[38][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane25_strm0_data          ( DownstreamStackBusLane[38][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane25_strm0_data_valid    ( DownstreamStackBusLane[38][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane25_strm1_ready         ( DownstreamStackBusLane[38][25].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane25_strm1_cntl          ( DownstreamStackBusLane[38][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane25_strm1_data          ( DownstreamStackBusLane[38][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane25_strm1_data_valid    ( DownstreamStackBusLane[38][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane26_strm0_ready         ( DownstreamStackBusLane[38][26].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane26_strm0_cntl          ( DownstreamStackBusLane[38][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane26_strm0_data          ( DownstreamStackBusLane[38][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane26_strm0_data_valid    ( DownstreamStackBusLane[38][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane26_strm1_ready         ( DownstreamStackBusLane[38][26].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane26_strm1_cntl          ( DownstreamStackBusLane[38][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane26_strm1_data          ( DownstreamStackBusLane[38][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane26_strm1_data_valid    ( DownstreamStackBusLane[38][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane27_strm0_ready         ( DownstreamStackBusLane[38][27].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane27_strm0_cntl          ( DownstreamStackBusLane[38][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane27_strm0_data          ( DownstreamStackBusLane[38][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane27_strm0_data_valid    ( DownstreamStackBusLane[38][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane27_strm1_ready         ( DownstreamStackBusLane[38][27].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane27_strm1_cntl          ( DownstreamStackBusLane[38][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane27_strm1_data          ( DownstreamStackBusLane[38][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane27_strm1_data_valid    ( DownstreamStackBusLane[38][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane28_strm0_ready         ( DownstreamStackBusLane[38][28].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane28_strm0_cntl          ( DownstreamStackBusLane[38][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane28_strm0_data          ( DownstreamStackBusLane[38][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane28_strm0_data_valid    ( DownstreamStackBusLane[38][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane28_strm1_ready         ( DownstreamStackBusLane[38][28].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane28_strm1_cntl          ( DownstreamStackBusLane[38][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane28_strm1_data          ( DownstreamStackBusLane[38][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane28_strm1_data_valid    ( DownstreamStackBusLane[38][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane29_strm0_ready         ( DownstreamStackBusLane[38][29].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane29_strm0_cntl          ( DownstreamStackBusLane[38][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane29_strm0_data          ( DownstreamStackBusLane[38][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane29_strm0_data_valid    ( DownstreamStackBusLane[38][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane29_strm1_ready         ( DownstreamStackBusLane[38][29].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane29_strm1_cntl          ( DownstreamStackBusLane[38][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane29_strm1_data          ( DownstreamStackBusLane[38][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane29_strm1_data_valid    ( DownstreamStackBusLane[38][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane30_strm0_ready         ( DownstreamStackBusLane[38][30].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane30_strm0_cntl          ( DownstreamStackBusLane[38][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane30_strm0_data          ( DownstreamStackBusLane[38][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane30_strm0_data_valid    ( DownstreamStackBusLane[38][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane30_strm1_ready         ( DownstreamStackBusLane[38][30].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane30_strm1_cntl          ( DownstreamStackBusLane[38][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane30_strm1_data          ( DownstreamStackBusLane[38][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane30_strm1_data_valid    ( DownstreamStackBusLane[38][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 38, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane31_strm0_ready         ( DownstreamStackBusLane[38][31].pe__std__lane_strm0_ready              ),      
        .std__pe38__lane31_strm0_cntl          ( DownstreamStackBusLane[38][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe38__lane31_strm0_data          ( DownstreamStackBusLane[38][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe38__lane31_strm0_data_valid    ( DownstreamStackBusLane[38][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__std__lane31_strm1_ready         ( DownstreamStackBusLane[38][31].pe__std__lane_strm1_ready              ),      
        .std__pe38__lane31_strm1_cntl          ( DownstreamStackBusLane[38][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe38__lane31_strm1_data          ( DownstreamStackBusLane[38][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe38__lane31_strm1_data_valid    ( DownstreamStackBusLane[38][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane0_strm0_ready         ( DownstreamStackBusLane[39][0].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane0_strm0_cntl          ( DownstreamStackBusLane[39][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane0_strm0_data          ( DownstreamStackBusLane[39][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane0_strm0_data_valid    ( DownstreamStackBusLane[39][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane0_strm1_ready         ( DownstreamStackBusLane[39][0].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane0_strm1_cntl          ( DownstreamStackBusLane[39][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane0_strm1_data          ( DownstreamStackBusLane[39][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane0_strm1_data_valid    ( DownstreamStackBusLane[39][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane1_strm0_ready         ( DownstreamStackBusLane[39][1].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane1_strm0_cntl          ( DownstreamStackBusLane[39][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane1_strm0_data          ( DownstreamStackBusLane[39][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane1_strm0_data_valid    ( DownstreamStackBusLane[39][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane1_strm1_ready         ( DownstreamStackBusLane[39][1].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane1_strm1_cntl          ( DownstreamStackBusLane[39][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane1_strm1_data          ( DownstreamStackBusLane[39][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane1_strm1_data_valid    ( DownstreamStackBusLane[39][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane2_strm0_ready         ( DownstreamStackBusLane[39][2].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane2_strm0_cntl          ( DownstreamStackBusLane[39][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane2_strm0_data          ( DownstreamStackBusLane[39][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane2_strm0_data_valid    ( DownstreamStackBusLane[39][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane2_strm1_ready         ( DownstreamStackBusLane[39][2].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane2_strm1_cntl          ( DownstreamStackBusLane[39][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane2_strm1_data          ( DownstreamStackBusLane[39][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane2_strm1_data_valid    ( DownstreamStackBusLane[39][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane3_strm0_ready         ( DownstreamStackBusLane[39][3].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane3_strm0_cntl          ( DownstreamStackBusLane[39][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane3_strm0_data          ( DownstreamStackBusLane[39][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane3_strm0_data_valid    ( DownstreamStackBusLane[39][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane3_strm1_ready         ( DownstreamStackBusLane[39][3].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane3_strm1_cntl          ( DownstreamStackBusLane[39][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane3_strm1_data          ( DownstreamStackBusLane[39][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane3_strm1_data_valid    ( DownstreamStackBusLane[39][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane4_strm0_ready         ( DownstreamStackBusLane[39][4].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane4_strm0_cntl          ( DownstreamStackBusLane[39][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane4_strm0_data          ( DownstreamStackBusLane[39][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane4_strm0_data_valid    ( DownstreamStackBusLane[39][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane4_strm1_ready         ( DownstreamStackBusLane[39][4].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane4_strm1_cntl          ( DownstreamStackBusLane[39][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane4_strm1_data          ( DownstreamStackBusLane[39][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane4_strm1_data_valid    ( DownstreamStackBusLane[39][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane5_strm0_ready         ( DownstreamStackBusLane[39][5].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane5_strm0_cntl          ( DownstreamStackBusLane[39][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane5_strm0_data          ( DownstreamStackBusLane[39][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane5_strm0_data_valid    ( DownstreamStackBusLane[39][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane5_strm1_ready         ( DownstreamStackBusLane[39][5].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane5_strm1_cntl          ( DownstreamStackBusLane[39][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane5_strm1_data          ( DownstreamStackBusLane[39][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane5_strm1_data_valid    ( DownstreamStackBusLane[39][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane6_strm0_ready         ( DownstreamStackBusLane[39][6].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane6_strm0_cntl          ( DownstreamStackBusLane[39][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane6_strm0_data          ( DownstreamStackBusLane[39][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane6_strm0_data_valid    ( DownstreamStackBusLane[39][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane6_strm1_ready         ( DownstreamStackBusLane[39][6].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane6_strm1_cntl          ( DownstreamStackBusLane[39][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane6_strm1_data          ( DownstreamStackBusLane[39][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane6_strm1_data_valid    ( DownstreamStackBusLane[39][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane7_strm0_ready         ( DownstreamStackBusLane[39][7].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane7_strm0_cntl          ( DownstreamStackBusLane[39][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane7_strm0_data          ( DownstreamStackBusLane[39][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane7_strm0_data_valid    ( DownstreamStackBusLane[39][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane7_strm1_ready         ( DownstreamStackBusLane[39][7].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane7_strm1_cntl          ( DownstreamStackBusLane[39][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane7_strm1_data          ( DownstreamStackBusLane[39][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane7_strm1_data_valid    ( DownstreamStackBusLane[39][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane8_strm0_ready         ( DownstreamStackBusLane[39][8].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane8_strm0_cntl          ( DownstreamStackBusLane[39][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane8_strm0_data          ( DownstreamStackBusLane[39][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane8_strm0_data_valid    ( DownstreamStackBusLane[39][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane8_strm1_ready         ( DownstreamStackBusLane[39][8].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane8_strm1_cntl          ( DownstreamStackBusLane[39][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane8_strm1_data          ( DownstreamStackBusLane[39][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane8_strm1_data_valid    ( DownstreamStackBusLane[39][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane9_strm0_ready         ( DownstreamStackBusLane[39][9].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane9_strm0_cntl          ( DownstreamStackBusLane[39][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane9_strm0_data          ( DownstreamStackBusLane[39][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane9_strm0_data_valid    ( DownstreamStackBusLane[39][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane9_strm1_ready         ( DownstreamStackBusLane[39][9].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane9_strm1_cntl          ( DownstreamStackBusLane[39][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane9_strm1_data          ( DownstreamStackBusLane[39][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane9_strm1_data_valid    ( DownstreamStackBusLane[39][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane10_strm0_ready         ( DownstreamStackBusLane[39][10].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane10_strm0_cntl          ( DownstreamStackBusLane[39][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane10_strm0_data          ( DownstreamStackBusLane[39][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane10_strm0_data_valid    ( DownstreamStackBusLane[39][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane10_strm1_ready         ( DownstreamStackBusLane[39][10].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane10_strm1_cntl          ( DownstreamStackBusLane[39][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane10_strm1_data          ( DownstreamStackBusLane[39][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane10_strm1_data_valid    ( DownstreamStackBusLane[39][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane11_strm0_ready         ( DownstreamStackBusLane[39][11].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane11_strm0_cntl          ( DownstreamStackBusLane[39][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane11_strm0_data          ( DownstreamStackBusLane[39][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane11_strm0_data_valid    ( DownstreamStackBusLane[39][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane11_strm1_ready         ( DownstreamStackBusLane[39][11].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane11_strm1_cntl          ( DownstreamStackBusLane[39][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane11_strm1_data          ( DownstreamStackBusLane[39][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane11_strm1_data_valid    ( DownstreamStackBusLane[39][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane12_strm0_ready         ( DownstreamStackBusLane[39][12].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane12_strm0_cntl          ( DownstreamStackBusLane[39][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane12_strm0_data          ( DownstreamStackBusLane[39][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane12_strm0_data_valid    ( DownstreamStackBusLane[39][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane12_strm1_ready         ( DownstreamStackBusLane[39][12].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane12_strm1_cntl          ( DownstreamStackBusLane[39][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane12_strm1_data          ( DownstreamStackBusLane[39][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane12_strm1_data_valid    ( DownstreamStackBusLane[39][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane13_strm0_ready         ( DownstreamStackBusLane[39][13].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane13_strm0_cntl          ( DownstreamStackBusLane[39][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane13_strm0_data          ( DownstreamStackBusLane[39][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane13_strm0_data_valid    ( DownstreamStackBusLane[39][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane13_strm1_ready         ( DownstreamStackBusLane[39][13].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane13_strm1_cntl          ( DownstreamStackBusLane[39][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane13_strm1_data          ( DownstreamStackBusLane[39][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane13_strm1_data_valid    ( DownstreamStackBusLane[39][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane14_strm0_ready         ( DownstreamStackBusLane[39][14].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane14_strm0_cntl          ( DownstreamStackBusLane[39][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane14_strm0_data          ( DownstreamStackBusLane[39][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane14_strm0_data_valid    ( DownstreamStackBusLane[39][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane14_strm1_ready         ( DownstreamStackBusLane[39][14].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane14_strm1_cntl          ( DownstreamStackBusLane[39][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane14_strm1_data          ( DownstreamStackBusLane[39][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane14_strm1_data_valid    ( DownstreamStackBusLane[39][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane15_strm0_ready         ( DownstreamStackBusLane[39][15].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane15_strm0_cntl          ( DownstreamStackBusLane[39][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane15_strm0_data          ( DownstreamStackBusLane[39][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane15_strm0_data_valid    ( DownstreamStackBusLane[39][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane15_strm1_ready         ( DownstreamStackBusLane[39][15].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane15_strm1_cntl          ( DownstreamStackBusLane[39][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane15_strm1_data          ( DownstreamStackBusLane[39][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane15_strm1_data_valid    ( DownstreamStackBusLane[39][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane16_strm0_ready         ( DownstreamStackBusLane[39][16].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane16_strm0_cntl          ( DownstreamStackBusLane[39][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane16_strm0_data          ( DownstreamStackBusLane[39][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane16_strm0_data_valid    ( DownstreamStackBusLane[39][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane16_strm1_ready         ( DownstreamStackBusLane[39][16].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane16_strm1_cntl          ( DownstreamStackBusLane[39][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane16_strm1_data          ( DownstreamStackBusLane[39][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane16_strm1_data_valid    ( DownstreamStackBusLane[39][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane17_strm0_ready         ( DownstreamStackBusLane[39][17].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane17_strm0_cntl          ( DownstreamStackBusLane[39][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane17_strm0_data          ( DownstreamStackBusLane[39][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane17_strm0_data_valid    ( DownstreamStackBusLane[39][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane17_strm1_ready         ( DownstreamStackBusLane[39][17].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane17_strm1_cntl          ( DownstreamStackBusLane[39][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane17_strm1_data          ( DownstreamStackBusLane[39][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane17_strm1_data_valid    ( DownstreamStackBusLane[39][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane18_strm0_ready         ( DownstreamStackBusLane[39][18].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane18_strm0_cntl          ( DownstreamStackBusLane[39][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane18_strm0_data          ( DownstreamStackBusLane[39][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane18_strm0_data_valid    ( DownstreamStackBusLane[39][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane18_strm1_ready         ( DownstreamStackBusLane[39][18].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane18_strm1_cntl          ( DownstreamStackBusLane[39][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane18_strm1_data          ( DownstreamStackBusLane[39][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane18_strm1_data_valid    ( DownstreamStackBusLane[39][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane19_strm0_ready         ( DownstreamStackBusLane[39][19].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane19_strm0_cntl          ( DownstreamStackBusLane[39][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane19_strm0_data          ( DownstreamStackBusLane[39][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane19_strm0_data_valid    ( DownstreamStackBusLane[39][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane19_strm1_ready         ( DownstreamStackBusLane[39][19].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane19_strm1_cntl          ( DownstreamStackBusLane[39][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane19_strm1_data          ( DownstreamStackBusLane[39][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane19_strm1_data_valid    ( DownstreamStackBusLane[39][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane20_strm0_ready         ( DownstreamStackBusLane[39][20].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane20_strm0_cntl          ( DownstreamStackBusLane[39][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane20_strm0_data          ( DownstreamStackBusLane[39][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane20_strm0_data_valid    ( DownstreamStackBusLane[39][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane20_strm1_ready         ( DownstreamStackBusLane[39][20].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane20_strm1_cntl          ( DownstreamStackBusLane[39][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane20_strm1_data          ( DownstreamStackBusLane[39][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane20_strm1_data_valid    ( DownstreamStackBusLane[39][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane21_strm0_ready         ( DownstreamStackBusLane[39][21].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane21_strm0_cntl          ( DownstreamStackBusLane[39][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane21_strm0_data          ( DownstreamStackBusLane[39][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane21_strm0_data_valid    ( DownstreamStackBusLane[39][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane21_strm1_ready         ( DownstreamStackBusLane[39][21].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane21_strm1_cntl          ( DownstreamStackBusLane[39][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane21_strm1_data          ( DownstreamStackBusLane[39][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane21_strm1_data_valid    ( DownstreamStackBusLane[39][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane22_strm0_ready         ( DownstreamStackBusLane[39][22].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane22_strm0_cntl          ( DownstreamStackBusLane[39][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane22_strm0_data          ( DownstreamStackBusLane[39][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane22_strm0_data_valid    ( DownstreamStackBusLane[39][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane22_strm1_ready         ( DownstreamStackBusLane[39][22].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane22_strm1_cntl          ( DownstreamStackBusLane[39][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane22_strm1_data          ( DownstreamStackBusLane[39][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane22_strm1_data_valid    ( DownstreamStackBusLane[39][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane23_strm0_ready         ( DownstreamStackBusLane[39][23].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane23_strm0_cntl          ( DownstreamStackBusLane[39][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane23_strm0_data          ( DownstreamStackBusLane[39][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane23_strm0_data_valid    ( DownstreamStackBusLane[39][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane23_strm1_ready         ( DownstreamStackBusLane[39][23].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane23_strm1_cntl          ( DownstreamStackBusLane[39][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane23_strm1_data          ( DownstreamStackBusLane[39][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane23_strm1_data_valid    ( DownstreamStackBusLane[39][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane24_strm0_ready         ( DownstreamStackBusLane[39][24].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane24_strm0_cntl          ( DownstreamStackBusLane[39][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane24_strm0_data          ( DownstreamStackBusLane[39][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane24_strm0_data_valid    ( DownstreamStackBusLane[39][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane24_strm1_ready         ( DownstreamStackBusLane[39][24].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane24_strm1_cntl          ( DownstreamStackBusLane[39][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane24_strm1_data          ( DownstreamStackBusLane[39][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane24_strm1_data_valid    ( DownstreamStackBusLane[39][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane25_strm0_ready         ( DownstreamStackBusLane[39][25].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane25_strm0_cntl          ( DownstreamStackBusLane[39][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane25_strm0_data          ( DownstreamStackBusLane[39][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane25_strm0_data_valid    ( DownstreamStackBusLane[39][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane25_strm1_ready         ( DownstreamStackBusLane[39][25].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane25_strm1_cntl          ( DownstreamStackBusLane[39][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane25_strm1_data          ( DownstreamStackBusLane[39][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane25_strm1_data_valid    ( DownstreamStackBusLane[39][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane26_strm0_ready         ( DownstreamStackBusLane[39][26].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane26_strm0_cntl          ( DownstreamStackBusLane[39][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane26_strm0_data          ( DownstreamStackBusLane[39][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane26_strm0_data_valid    ( DownstreamStackBusLane[39][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane26_strm1_ready         ( DownstreamStackBusLane[39][26].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane26_strm1_cntl          ( DownstreamStackBusLane[39][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane26_strm1_data          ( DownstreamStackBusLane[39][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane26_strm1_data_valid    ( DownstreamStackBusLane[39][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane27_strm0_ready         ( DownstreamStackBusLane[39][27].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane27_strm0_cntl          ( DownstreamStackBusLane[39][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane27_strm0_data          ( DownstreamStackBusLane[39][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane27_strm0_data_valid    ( DownstreamStackBusLane[39][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane27_strm1_ready         ( DownstreamStackBusLane[39][27].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane27_strm1_cntl          ( DownstreamStackBusLane[39][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane27_strm1_data          ( DownstreamStackBusLane[39][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane27_strm1_data_valid    ( DownstreamStackBusLane[39][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane28_strm0_ready         ( DownstreamStackBusLane[39][28].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane28_strm0_cntl          ( DownstreamStackBusLane[39][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane28_strm0_data          ( DownstreamStackBusLane[39][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane28_strm0_data_valid    ( DownstreamStackBusLane[39][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane28_strm1_ready         ( DownstreamStackBusLane[39][28].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane28_strm1_cntl          ( DownstreamStackBusLane[39][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane28_strm1_data          ( DownstreamStackBusLane[39][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane28_strm1_data_valid    ( DownstreamStackBusLane[39][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane29_strm0_ready         ( DownstreamStackBusLane[39][29].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane29_strm0_cntl          ( DownstreamStackBusLane[39][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane29_strm0_data          ( DownstreamStackBusLane[39][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane29_strm0_data_valid    ( DownstreamStackBusLane[39][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane29_strm1_ready         ( DownstreamStackBusLane[39][29].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane29_strm1_cntl          ( DownstreamStackBusLane[39][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane29_strm1_data          ( DownstreamStackBusLane[39][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane29_strm1_data_valid    ( DownstreamStackBusLane[39][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane30_strm0_ready         ( DownstreamStackBusLane[39][30].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane30_strm0_cntl          ( DownstreamStackBusLane[39][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane30_strm0_data          ( DownstreamStackBusLane[39][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane30_strm0_data_valid    ( DownstreamStackBusLane[39][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane30_strm1_ready         ( DownstreamStackBusLane[39][30].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane30_strm1_cntl          ( DownstreamStackBusLane[39][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane30_strm1_data          ( DownstreamStackBusLane[39][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane30_strm1_data_valid    ( DownstreamStackBusLane[39][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 39, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane31_strm0_ready         ( DownstreamStackBusLane[39][31].pe__std__lane_strm0_ready              ),      
        .std__pe39__lane31_strm0_cntl          ( DownstreamStackBusLane[39][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe39__lane31_strm0_data          ( DownstreamStackBusLane[39][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe39__lane31_strm0_data_valid    ( DownstreamStackBusLane[39][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__std__lane31_strm1_ready         ( DownstreamStackBusLane[39][31].pe__std__lane_strm1_ready              ),      
        .std__pe39__lane31_strm1_cntl          ( DownstreamStackBusLane[39][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe39__lane31_strm1_data          ( DownstreamStackBusLane[39][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe39__lane31_strm1_data_valid    ( DownstreamStackBusLane[39][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane0_strm0_ready         ( DownstreamStackBusLane[40][0].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane0_strm0_cntl          ( DownstreamStackBusLane[40][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane0_strm0_data          ( DownstreamStackBusLane[40][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane0_strm0_data_valid    ( DownstreamStackBusLane[40][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane0_strm1_ready         ( DownstreamStackBusLane[40][0].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane0_strm1_cntl          ( DownstreamStackBusLane[40][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane0_strm1_data          ( DownstreamStackBusLane[40][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane0_strm1_data_valid    ( DownstreamStackBusLane[40][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane1_strm0_ready         ( DownstreamStackBusLane[40][1].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane1_strm0_cntl          ( DownstreamStackBusLane[40][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane1_strm0_data          ( DownstreamStackBusLane[40][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane1_strm0_data_valid    ( DownstreamStackBusLane[40][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane1_strm1_ready         ( DownstreamStackBusLane[40][1].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane1_strm1_cntl          ( DownstreamStackBusLane[40][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane1_strm1_data          ( DownstreamStackBusLane[40][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane1_strm1_data_valid    ( DownstreamStackBusLane[40][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane2_strm0_ready         ( DownstreamStackBusLane[40][2].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane2_strm0_cntl          ( DownstreamStackBusLane[40][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane2_strm0_data          ( DownstreamStackBusLane[40][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane2_strm0_data_valid    ( DownstreamStackBusLane[40][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane2_strm1_ready         ( DownstreamStackBusLane[40][2].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane2_strm1_cntl          ( DownstreamStackBusLane[40][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane2_strm1_data          ( DownstreamStackBusLane[40][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane2_strm1_data_valid    ( DownstreamStackBusLane[40][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane3_strm0_ready         ( DownstreamStackBusLane[40][3].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane3_strm0_cntl          ( DownstreamStackBusLane[40][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane3_strm0_data          ( DownstreamStackBusLane[40][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane3_strm0_data_valid    ( DownstreamStackBusLane[40][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane3_strm1_ready         ( DownstreamStackBusLane[40][3].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane3_strm1_cntl          ( DownstreamStackBusLane[40][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane3_strm1_data          ( DownstreamStackBusLane[40][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane3_strm1_data_valid    ( DownstreamStackBusLane[40][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane4_strm0_ready         ( DownstreamStackBusLane[40][4].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane4_strm0_cntl          ( DownstreamStackBusLane[40][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane4_strm0_data          ( DownstreamStackBusLane[40][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane4_strm0_data_valid    ( DownstreamStackBusLane[40][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane4_strm1_ready         ( DownstreamStackBusLane[40][4].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane4_strm1_cntl          ( DownstreamStackBusLane[40][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane4_strm1_data          ( DownstreamStackBusLane[40][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane4_strm1_data_valid    ( DownstreamStackBusLane[40][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane5_strm0_ready         ( DownstreamStackBusLane[40][5].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane5_strm0_cntl          ( DownstreamStackBusLane[40][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane5_strm0_data          ( DownstreamStackBusLane[40][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane5_strm0_data_valid    ( DownstreamStackBusLane[40][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane5_strm1_ready         ( DownstreamStackBusLane[40][5].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane5_strm1_cntl          ( DownstreamStackBusLane[40][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane5_strm1_data          ( DownstreamStackBusLane[40][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane5_strm1_data_valid    ( DownstreamStackBusLane[40][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane6_strm0_ready         ( DownstreamStackBusLane[40][6].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane6_strm0_cntl          ( DownstreamStackBusLane[40][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane6_strm0_data          ( DownstreamStackBusLane[40][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane6_strm0_data_valid    ( DownstreamStackBusLane[40][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane6_strm1_ready         ( DownstreamStackBusLane[40][6].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane6_strm1_cntl          ( DownstreamStackBusLane[40][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane6_strm1_data          ( DownstreamStackBusLane[40][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane6_strm1_data_valid    ( DownstreamStackBusLane[40][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane7_strm0_ready         ( DownstreamStackBusLane[40][7].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane7_strm0_cntl          ( DownstreamStackBusLane[40][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane7_strm0_data          ( DownstreamStackBusLane[40][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane7_strm0_data_valid    ( DownstreamStackBusLane[40][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane7_strm1_ready         ( DownstreamStackBusLane[40][7].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane7_strm1_cntl          ( DownstreamStackBusLane[40][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane7_strm1_data          ( DownstreamStackBusLane[40][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane7_strm1_data_valid    ( DownstreamStackBusLane[40][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane8_strm0_ready         ( DownstreamStackBusLane[40][8].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane8_strm0_cntl          ( DownstreamStackBusLane[40][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane8_strm0_data          ( DownstreamStackBusLane[40][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane8_strm0_data_valid    ( DownstreamStackBusLane[40][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane8_strm1_ready         ( DownstreamStackBusLane[40][8].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane8_strm1_cntl          ( DownstreamStackBusLane[40][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane8_strm1_data          ( DownstreamStackBusLane[40][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane8_strm1_data_valid    ( DownstreamStackBusLane[40][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane9_strm0_ready         ( DownstreamStackBusLane[40][9].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane9_strm0_cntl          ( DownstreamStackBusLane[40][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane9_strm0_data          ( DownstreamStackBusLane[40][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane9_strm0_data_valid    ( DownstreamStackBusLane[40][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane9_strm1_ready         ( DownstreamStackBusLane[40][9].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane9_strm1_cntl          ( DownstreamStackBusLane[40][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane9_strm1_data          ( DownstreamStackBusLane[40][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane9_strm1_data_valid    ( DownstreamStackBusLane[40][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane10_strm0_ready         ( DownstreamStackBusLane[40][10].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane10_strm0_cntl          ( DownstreamStackBusLane[40][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane10_strm0_data          ( DownstreamStackBusLane[40][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane10_strm0_data_valid    ( DownstreamStackBusLane[40][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane10_strm1_ready         ( DownstreamStackBusLane[40][10].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane10_strm1_cntl          ( DownstreamStackBusLane[40][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane10_strm1_data          ( DownstreamStackBusLane[40][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane10_strm1_data_valid    ( DownstreamStackBusLane[40][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane11_strm0_ready         ( DownstreamStackBusLane[40][11].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane11_strm0_cntl          ( DownstreamStackBusLane[40][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane11_strm0_data          ( DownstreamStackBusLane[40][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane11_strm0_data_valid    ( DownstreamStackBusLane[40][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane11_strm1_ready         ( DownstreamStackBusLane[40][11].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane11_strm1_cntl          ( DownstreamStackBusLane[40][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane11_strm1_data          ( DownstreamStackBusLane[40][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane11_strm1_data_valid    ( DownstreamStackBusLane[40][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane12_strm0_ready         ( DownstreamStackBusLane[40][12].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane12_strm0_cntl          ( DownstreamStackBusLane[40][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane12_strm0_data          ( DownstreamStackBusLane[40][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane12_strm0_data_valid    ( DownstreamStackBusLane[40][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane12_strm1_ready         ( DownstreamStackBusLane[40][12].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane12_strm1_cntl          ( DownstreamStackBusLane[40][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane12_strm1_data          ( DownstreamStackBusLane[40][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane12_strm1_data_valid    ( DownstreamStackBusLane[40][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane13_strm0_ready         ( DownstreamStackBusLane[40][13].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane13_strm0_cntl          ( DownstreamStackBusLane[40][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane13_strm0_data          ( DownstreamStackBusLane[40][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane13_strm0_data_valid    ( DownstreamStackBusLane[40][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane13_strm1_ready         ( DownstreamStackBusLane[40][13].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane13_strm1_cntl          ( DownstreamStackBusLane[40][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane13_strm1_data          ( DownstreamStackBusLane[40][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane13_strm1_data_valid    ( DownstreamStackBusLane[40][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane14_strm0_ready         ( DownstreamStackBusLane[40][14].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane14_strm0_cntl          ( DownstreamStackBusLane[40][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane14_strm0_data          ( DownstreamStackBusLane[40][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane14_strm0_data_valid    ( DownstreamStackBusLane[40][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane14_strm1_ready         ( DownstreamStackBusLane[40][14].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane14_strm1_cntl          ( DownstreamStackBusLane[40][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane14_strm1_data          ( DownstreamStackBusLane[40][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane14_strm1_data_valid    ( DownstreamStackBusLane[40][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane15_strm0_ready         ( DownstreamStackBusLane[40][15].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane15_strm0_cntl          ( DownstreamStackBusLane[40][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane15_strm0_data          ( DownstreamStackBusLane[40][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane15_strm0_data_valid    ( DownstreamStackBusLane[40][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane15_strm1_ready         ( DownstreamStackBusLane[40][15].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane15_strm1_cntl          ( DownstreamStackBusLane[40][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane15_strm1_data          ( DownstreamStackBusLane[40][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane15_strm1_data_valid    ( DownstreamStackBusLane[40][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane16_strm0_ready         ( DownstreamStackBusLane[40][16].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane16_strm0_cntl          ( DownstreamStackBusLane[40][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane16_strm0_data          ( DownstreamStackBusLane[40][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane16_strm0_data_valid    ( DownstreamStackBusLane[40][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane16_strm1_ready         ( DownstreamStackBusLane[40][16].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane16_strm1_cntl          ( DownstreamStackBusLane[40][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane16_strm1_data          ( DownstreamStackBusLane[40][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane16_strm1_data_valid    ( DownstreamStackBusLane[40][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane17_strm0_ready         ( DownstreamStackBusLane[40][17].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane17_strm0_cntl          ( DownstreamStackBusLane[40][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane17_strm0_data          ( DownstreamStackBusLane[40][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane17_strm0_data_valid    ( DownstreamStackBusLane[40][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane17_strm1_ready         ( DownstreamStackBusLane[40][17].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane17_strm1_cntl          ( DownstreamStackBusLane[40][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane17_strm1_data          ( DownstreamStackBusLane[40][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane17_strm1_data_valid    ( DownstreamStackBusLane[40][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane18_strm0_ready         ( DownstreamStackBusLane[40][18].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane18_strm0_cntl          ( DownstreamStackBusLane[40][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane18_strm0_data          ( DownstreamStackBusLane[40][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane18_strm0_data_valid    ( DownstreamStackBusLane[40][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane18_strm1_ready         ( DownstreamStackBusLane[40][18].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane18_strm1_cntl          ( DownstreamStackBusLane[40][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane18_strm1_data          ( DownstreamStackBusLane[40][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane18_strm1_data_valid    ( DownstreamStackBusLane[40][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane19_strm0_ready         ( DownstreamStackBusLane[40][19].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane19_strm0_cntl          ( DownstreamStackBusLane[40][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane19_strm0_data          ( DownstreamStackBusLane[40][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane19_strm0_data_valid    ( DownstreamStackBusLane[40][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane19_strm1_ready         ( DownstreamStackBusLane[40][19].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane19_strm1_cntl          ( DownstreamStackBusLane[40][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane19_strm1_data          ( DownstreamStackBusLane[40][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane19_strm1_data_valid    ( DownstreamStackBusLane[40][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane20_strm0_ready         ( DownstreamStackBusLane[40][20].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane20_strm0_cntl          ( DownstreamStackBusLane[40][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane20_strm0_data          ( DownstreamStackBusLane[40][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane20_strm0_data_valid    ( DownstreamStackBusLane[40][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane20_strm1_ready         ( DownstreamStackBusLane[40][20].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane20_strm1_cntl          ( DownstreamStackBusLane[40][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane20_strm1_data          ( DownstreamStackBusLane[40][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane20_strm1_data_valid    ( DownstreamStackBusLane[40][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane21_strm0_ready         ( DownstreamStackBusLane[40][21].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane21_strm0_cntl          ( DownstreamStackBusLane[40][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane21_strm0_data          ( DownstreamStackBusLane[40][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane21_strm0_data_valid    ( DownstreamStackBusLane[40][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane21_strm1_ready         ( DownstreamStackBusLane[40][21].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane21_strm1_cntl          ( DownstreamStackBusLane[40][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane21_strm1_data          ( DownstreamStackBusLane[40][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane21_strm1_data_valid    ( DownstreamStackBusLane[40][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane22_strm0_ready         ( DownstreamStackBusLane[40][22].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane22_strm0_cntl          ( DownstreamStackBusLane[40][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane22_strm0_data          ( DownstreamStackBusLane[40][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane22_strm0_data_valid    ( DownstreamStackBusLane[40][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane22_strm1_ready         ( DownstreamStackBusLane[40][22].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane22_strm1_cntl          ( DownstreamStackBusLane[40][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane22_strm1_data          ( DownstreamStackBusLane[40][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane22_strm1_data_valid    ( DownstreamStackBusLane[40][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane23_strm0_ready         ( DownstreamStackBusLane[40][23].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane23_strm0_cntl          ( DownstreamStackBusLane[40][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane23_strm0_data          ( DownstreamStackBusLane[40][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane23_strm0_data_valid    ( DownstreamStackBusLane[40][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane23_strm1_ready         ( DownstreamStackBusLane[40][23].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane23_strm1_cntl          ( DownstreamStackBusLane[40][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane23_strm1_data          ( DownstreamStackBusLane[40][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane23_strm1_data_valid    ( DownstreamStackBusLane[40][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane24_strm0_ready         ( DownstreamStackBusLane[40][24].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane24_strm0_cntl          ( DownstreamStackBusLane[40][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane24_strm0_data          ( DownstreamStackBusLane[40][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane24_strm0_data_valid    ( DownstreamStackBusLane[40][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane24_strm1_ready         ( DownstreamStackBusLane[40][24].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane24_strm1_cntl          ( DownstreamStackBusLane[40][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane24_strm1_data          ( DownstreamStackBusLane[40][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane24_strm1_data_valid    ( DownstreamStackBusLane[40][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane25_strm0_ready         ( DownstreamStackBusLane[40][25].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane25_strm0_cntl          ( DownstreamStackBusLane[40][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane25_strm0_data          ( DownstreamStackBusLane[40][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane25_strm0_data_valid    ( DownstreamStackBusLane[40][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane25_strm1_ready         ( DownstreamStackBusLane[40][25].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane25_strm1_cntl          ( DownstreamStackBusLane[40][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane25_strm1_data          ( DownstreamStackBusLane[40][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane25_strm1_data_valid    ( DownstreamStackBusLane[40][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane26_strm0_ready         ( DownstreamStackBusLane[40][26].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane26_strm0_cntl          ( DownstreamStackBusLane[40][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane26_strm0_data          ( DownstreamStackBusLane[40][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane26_strm0_data_valid    ( DownstreamStackBusLane[40][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane26_strm1_ready         ( DownstreamStackBusLane[40][26].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane26_strm1_cntl          ( DownstreamStackBusLane[40][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane26_strm1_data          ( DownstreamStackBusLane[40][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane26_strm1_data_valid    ( DownstreamStackBusLane[40][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane27_strm0_ready         ( DownstreamStackBusLane[40][27].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane27_strm0_cntl          ( DownstreamStackBusLane[40][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane27_strm0_data          ( DownstreamStackBusLane[40][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane27_strm0_data_valid    ( DownstreamStackBusLane[40][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane27_strm1_ready         ( DownstreamStackBusLane[40][27].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane27_strm1_cntl          ( DownstreamStackBusLane[40][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane27_strm1_data          ( DownstreamStackBusLane[40][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane27_strm1_data_valid    ( DownstreamStackBusLane[40][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane28_strm0_ready         ( DownstreamStackBusLane[40][28].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane28_strm0_cntl          ( DownstreamStackBusLane[40][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane28_strm0_data          ( DownstreamStackBusLane[40][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane28_strm0_data_valid    ( DownstreamStackBusLane[40][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane28_strm1_ready         ( DownstreamStackBusLane[40][28].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane28_strm1_cntl          ( DownstreamStackBusLane[40][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane28_strm1_data          ( DownstreamStackBusLane[40][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane28_strm1_data_valid    ( DownstreamStackBusLane[40][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane29_strm0_ready         ( DownstreamStackBusLane[40][29].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane29_strm0_cntl          ( DownstreamStackBusLane[40][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane29_strm0_data          ( DownstreamStackBusLane[40][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane29_strm0_data_valid    ( DownstreamStackBusLane[40][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane29_strm1_ready         ( DownstreamStackBusLane[40][29].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane29_strm1_cntl          ( DownstreamStackBusLane[40][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane29_strm1_data          ( DownstreamStackBusLane[40][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane29_strm1_data_valid    ( DownstreamStackBusLane[40][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane30_strm0_ready         ( DownstreamStackBusLane[40][30].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane30_strm0_cntl          ( DownstreamStackBusLane[40][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane30_strm0_data          ( DownstreamStackBusLane[40][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane30_strm0_data_valid    ( DownstreamStackBusLane[40][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane30_strm1_ready         ( DownstreamStackBusLane[40][30].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane30_strm1_cntl          ( DownstreamStackBusLane[40][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane30_strm1_data          ( DownstreamStackBusLane[40][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane30_strm1_data_valid    ( DownstreamStackBusLane[40][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 40, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane31_strm0_ready         ( DownstreamStackBusLane[40][31].pe__std__lane_strm0_ready              ),      
        .std__pe40__lane31_strm0_cntl          ( DownstreamStackBusLane[40][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe40__lane31_strm0_data          ( DownstreamStackBusLane[40][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe40__lane31_strm0_data_valid    ( DownstreamStackBusLane[40][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__std__lane31_strm1_ready         ( DownstreamStackBusLane[40][31].pe__std__lane_strm1_ready              ),      
        .std__pe40__lane31_strm1_cntl          ( DownstreamStackBusLane[40][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe40__lane31_strm1_data          ( DownstreamStackBusLane[40][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe40__lane31_strm1_data_valid    ( DownstreamStackBusLane[40][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane0_strm0_ready         ( DownstreamStackBusLane[41][0].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane0_strm0_cntl          ( DownstreamStackBusLane[41][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane0_strm0_data          ( DownstreamStackBusLane[41][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane0_strm0_data_valid    ( DownstreamStackBusLane[41][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane0_strm1_ready         ( DownstreamStackBusLane[41][0].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane0_strm1_cntl          ( DownstreamStackBusLane[41][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane0_strm1_data          ( DownstreamStackBusLane[41][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane0_strm1_data_valid    ( DownstreamStackBusLane[41][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane1_strm0_ready         ( DownstreamStackBusLane[41][1].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane1_strm0_cntl          ( DownstreamStackBusLane[41][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane1_strm0_data          ( DownstreamStackBusLane[41][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane1_strm0_data_valid    ( DownstreamStackBusLane[41][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane1_strm1_ready         ( DownstreamStackBusLane[41][1].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane1_strm1_cntl          ( DownstreamStackBusLane[41][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane1_strm1_data          ( DownstreamStackBusLane[41][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane1_strm1_data_valid    ( DownstreamStackBusLane[41][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane2_strm0_ready         ( DownstreamStackBusLane[41][2].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane2_strm0_cntl          ( DownstreamStackBusLane[41][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane2_strm0_data          ( DownstreamStackBusLane[41][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane2_strm0_data_valid    ( DownstreamStackBusLane[41][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane2_strm1_ready         ( DownstreamStackBusLane[41][2].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane2_strm1_cntl          ( DownstreamStackBusLane[41][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane2_strm1_data          ( DownstreamStackBusLane[41][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane2_strm1_data_valid    ( DownstreamStackBusLane[41][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane3_strm0_ready         ( DownstreamStackBusLane[41][3].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane3_strm0_cntl          ( DownstreamStackBusLane[41][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane3_strm0_data          ( DownstreamStackBusLane[41][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane3_strm0_data_valid    ( DownstreamStackBusLane[41][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane3_strm1_ready         ( DownstreamStackBusLane[41][3].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane3_strm1_cntl          ( DownstreamStackBusLane[41][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane3_strm1_data          ( DownstreamStackBusLane[41][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane3_strm1_data_valid    ( DownstreamStackBusLane[41][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane4_strm0_ready         ( DownstreamStackBusLane[41][4].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane4_strm0_cntl          ( DownstreamStackBusLane[41][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane4_strm0_data          ( DownstreamStackBusLane[41][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane4_strm0_data_valid    ( DownstreamStackBusLane[41][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane4_strm1_ready         ( DownstreamStackBusLane[41][4].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane4_strm1_cntl          ( DownstreamStackBusLane[41][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane4_strm1_data          ( DownstreamStackBusLane[41][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane4_strm1_data_valid    ( DownstreamStackBusLane[41][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane5_strm0_ready         ( DownstreamStackBusLane[41][5].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane5_strm0_cntl          ( DownstreamStackBusLane[41][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane5_strm0_data          ( DownstreamStackBusLane[41][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane5_strm0_data_valid    ( DownstreamStackBusLane[41][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane5_strm1_ready         ( DownstreamStackBusLane[41][5].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane5_strm1_cntl          ( DownstreamStackBusLane[41][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane5_strm1_data          ( DownstreamStackBusLane[41][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane5_strm1_data_valid    ( DownstreamStackBusLane[41][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane6_strm0_ready         ( DownstreamStackBusLane[41][6].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane6_strm0_cntl          ( DownstreamStackBusLane[41][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane6_strm0_data          ( DownstreamStackBusLane[41][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane6_strm0_data_valid    ( DownstreamStackBusLane[41][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane6_strm1_ready         ( DownstreamStackBusLane[41][6].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane6_strm1_cntl          ( DownstreamStackBusLane[41][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane6_strm1_data          ( DownstreamStackBusLane[41][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane6_strm1_data_valid    ( DownstreamStackBusLane[41][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane7_strm0_ready         ( DownstreamStackBusLane[41][7].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane7_strm0_cntl          ( DownstreamStackBusLane[41][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane7_strm0_data          ( DownstreamStackBusLane[41][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane7_strm0_data_valid    ( DownstreamStackBusLane[41][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane7_strm1_ready         ( DownstreamStackBusLane[41][7].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane7_strm1_cntl          ( DownstreamStackBusLane[41][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane7_strm1_data          ( DownstreamStackBusLane[41][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane7_strm1_data_valid    ( DownstreamStackBusLane[41][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane8_strm0_ready         ( DownstreamStackBusLane[41][8].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane8_strm0_cntl          ( DownstreamStackBusLane[41][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane8_strm0_data          ( DownstreamStackBusLane[41][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane8_strm0_data_valid    ( DownstreamStackBusLane[41][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane8_strm1_ready         ( DownstreamStackBusLane[41][8].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane8_strm1_cntl          ( DownstreamStackBusLane[41][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane8_strm1_data          ( DownstreamStackBusLane[41][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane8_strm1_data_valid    ( DownstreamStackBusLane[41][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane9_strm0_ready         ( DownstreamStackBusLane[41][9].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane9_strm0_cntl          ( DownstreamStackBusLane[41][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane9_strm0_data          ( DownstreamStackBusLane[41][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane9_strm0_data_valid    ( DownstreamStackBusLane[41][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane9_strm1_ready         ( DownstreamStackBusLane[41][9].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane9_strm1_cntl          ( DownstreamStackBusLane[41][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane9_strm1_data          ( DownstreamStackBusLane[41][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane9_strm1_data_valid    ( DownstreamStackBusLane[41][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane10_strm0_ready         ( DownstreamStackBusLane[41][10].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane10_strm0_cntl          ( DownstreamStackBusLane[41][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane10_strm0_data          ( DownstreamStackBusLane[41][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane10_strm0_data_valid    ( DownstreamStackBusLane[41][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane10_strm1_ready         ( DownstreamStackBusLane[41][10].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane10_strm1_cntl          ( DownstreamStackBusLane[41][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane10_strm1_data          ( DownstreamStackBusLane[41][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane10_strm1_data_valid    ( DownstreamStackBusLane[41][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane11_strm0_ready         ( DownstreamStackBusLane[41][11].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane11_strm0_cntl          ( DownstreamStackBusLane[41][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane11_strm0_data          ( DownstreamStackBusLane[41][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane11_strm0_data_valid    ( DownstreamStackBusLane[41][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane11_strm1_ready         ( DownstreamStackBusLane[41][11].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane11_strm1_cntl          ( DownstreamStackBusLane[41][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane11_strm1_data          ( DownstreamStackBusLane[41][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane11_strm1_data_valid    ( DownstreamStackBusLane[41][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane12_strm0_ready         ( DownstreamStackBusLane[41][12].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane12_strm0_cntl          ( DownstreamStackBusLane[41][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane12_strm0_data          ( DownstreamStackBusLane[41][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane12_strm0_data_valid    ( DownstreamStackBusLane[41][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane12_strm1_ready         ( DownstreamStackBusLane[41][12].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane12_strm1_cntl          ( DownstreamStackBusLane[41][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane12_strm1_data          ( DownstreamStackBusLane[41][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane12_strm1_data_valid    ( DownstreamStackBusLane[41][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane13_strm0_ready         ( DownstreamStackBusLane[41][13].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane13_strm0_cntl          ( DownstreamStackBusLane[41][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane13_strm0_data          ( DownstreamStackBusLane[41][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane13_strm0_data_valid    ( DownstreamStackBusLane[41][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane13_strm1_ready         ( DownstreamStackBusLane[41][13].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane13_strm1_cntl          ( DownstreamStackBusLane[41][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane13_strm1_data          ( DownstreamStackBusLane[41][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane13_strm1_data_valid    ( DownstreamStackBusLane[41][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane14_strm0_ready         ( DownstreamStackBusLane[41][14].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane14_strm0_cntl          ( DownstreamStackBusLane[41][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane14_strm0_data          ( DownstreamStackBusLane[41][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane14_strm0_data_valid    ( DownstreamStackBusLane[41][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane14_strm1_ready         ( DownstreamStackBusLane[41][14].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane14_strm1_cntl          ( DownstreamStackBusLane[41][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane14_strm1_data          ( DownstreamStackBusLane[41][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane14_strm1_data_valid    ( DownstreamStackBusLane[41][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane15_strm0_ready         ( DownstreamStackBusLane[41][15].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane15_strm0_cntl          ( DownstreamStackBusLane[41][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane15_strm0_data          ( DownstreamStackBusLane[41][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane15_strm0_data_valid    ( DownstreamStackBusLane[41][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane15_strm1_ready         ( DownstreamStackBusLane[41][15].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane15_strm1_cntl          ( DownstreamStackBusLane[41][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane15_strm1_data          ( DownstreamStackBusLane[41][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane15_strm1_data_valid    ( DownstreamStackBusLane[41][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane16_strm0_ready         ( DownstreamStackBusLane[41][16].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane16_strm0_cntl          ( DownstreamStackBusLane[41][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane16_strm0_data          ( DownstreamStackBusLane[41][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane16_strm0_data_valid    ( DownstreamStackBusLane[41][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane16_strm1_ready         ( DownstreamStackBusLane[41][16].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane16_strm1_cntl          ( DownstreamStackBusLane[41][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane16_strm1_data          ( DownstreamStackBusLane[41][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane16_strm1_data_valid    ( DownstreamStackBusLane[41][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane17_strm0_ready         ( DownstreamStackBusLane[41][17].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane17_strm0_cntl          ( DownstreamStackBusLane[41][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane17_strm0_data          ( DownstreamStackBusLane[41][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane17_strm0_data_valid    ( DownstreamStackBusLane[41][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane17_strm1_ready         ( DownstreamStackBusLane[41][17].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane17_strm1_cntl          ( DownstreamStackBusLane[41][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane17_strm1_data          ( DownstreamStackBusLane[41][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane17_strm1_data_valid    ( DownstreamStackBusLane[41][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane18_strm0_ready         ( DownstreamStackBusLane[41][18].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane18_strm0_cntl          ( DownstreamStackBusLane[41][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane18_strm0_data          ( DownstreamStackBusLane[41][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane18_strm0_data_valid    ( DownstreamStackBusLane[41][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane18_strm1_ready         ( DownstreamStackBusLane[41][18].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane18_strm1_cntl          ( DownstreamStackBusLane[41][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane18_strm1_data          ( DownstreamStackBusLane[41][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane18_strm1_data_valid    ( DownstreamStackBusLane[41][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane19_strm0_ready         ( DownstreamStackBusLane[41][19].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane19_strm0_cntl          ( DownstreamStackBusLane[41][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane19_strm0_data          ( DownstreamStackBusLane[41][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane19_strm0_data_valid    ( DownstreamStackBusLane[41][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane19_strm1_ready         ( DownstreamStackBusLane[41][19].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane19_strm1_cntl          ( DownstreamStackBusLane[41][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane19_strm1_data          ( DownstreamStackBusLane[41][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane19_strm1_data_valid    ( DownstreamStackBusLane[41][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane20_strm0_ready         ( DownstreamStackBusLane[41][20].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane20_strm0_cntl          ( DownstreamStackBusLane[41][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane20_strm0_data          ( DownstreamStackBusLane[41][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane20_strm0_data_valid    ( DownstreamStackBusLane[41][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane20_strm1_ready         ( DownstreamStackBusLane[41][20].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane20_strm1_cntl          ( DownstreamStackBusLane[41][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane20_strm1_data          ( DownstreamStackBusLane[41][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane20_strm1_data_valid    ( DownstreamStackBusLane[41][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane21_strm0_ready         ( DownstreamStackBusLane[41][21].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane21_strm0_cntl          ( DownstreamStackBusLane[41][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane21_strm0_data          ( DownstreamStackBusLane[41][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane21_strm0_data_valid    ( DownstreamStackBusLane[41][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane21_strm1_ready         ( DownstreamStackBusLane[41][21].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane21_strm1_cntl          ( DownstreamStackBusLane[41][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane21_strm1_data          ( DownstreamStackBusLane[41][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane21_strm1_data_valid    ( DownstreamStackBusLane[41][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane22_strm0_ready         ( DownstreamStackBusLane[41][22].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane22_strm0_cntl          ( DownstreamStackBusLane[41][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane22_strm0_data          ( DownstreamStackBusLane[41][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane22_strm0_data_valid    ( DownstreamStackBusLane[41][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane22_strm1_ready         ( DownstreamStackBusLane[41][22].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane22_strm1_cntl          ( DownstreamStackBusLane[41][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane22_strm1_data          ( DownstreamStackBusLane[41][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane22_strm1_data_valid    ( DownstreamStackBusLane[41][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane23_strm0_ready         ( DownstreamStackBusLane[41][23].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane23_strm0_cntl          ( DownstreamStackBusLane[41][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane23_strm0_data          ( DownstreamStackBusLane[41][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane23_strm0_data_valid    ( DownstreamStackBusLane[41][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane23_strm1_ready         ( DownstreamStackBusLane[41][23].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane23_strm1_cntl          ( DownstreamStackBusLane[41][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane23_strm1_data          ( DownstreamStackBusLane[41][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane23_strm1_data_valid    ( DownstreamStackBusLane[41][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane24_strm0_ready         ( DownstreamStackBusLane[41][24].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane24_strm0_cntl          ( DownstreamStackBusLane[41][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane24_strm0_data          ( DownstreamStackBusLane[41][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane24_strm0_data_valid    ( DownstreamStackBusLane[41][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane24_strm1_ready         ( DownstreamStackBusLane[41][24].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane24_strm1_cntl          ( DownstreamStackBusLane[41][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane24_strm1_data          ( DownstreamStackBusLane[41][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane24_strm1_data_valid    ( DownstreamStackBusLane[41][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane25_strm0_ready         ( DownstreamStackBusLane[41][25].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane25_strm0_cntl          ( DownstreamStackBusLane[41][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane25_strm0_data          ( DownstreamStackBusLane[41][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane25_strm0_data_valid    ( DownstreamStackBusLane[41][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane25_strm1_ready         ( DownstreamStackBusLane[41][25].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane25_strm1_cntl          ( DownstreamStackBusLane[41][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane25_strm1_data          ( DownstreamStackBusLane[41][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane25_strm1_data_valid    ( DownstreamStackBusLane[41][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane26_strm0_ready         ( DownstreamStackBusLane[41][26].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane26_strm0_cntl          ( DownstreamStackBusLane[41][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane26_strm0_data          ( DownstreamStackBusLane[41][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane26_strm0_data_valid    ( DownstreamStackBusLane[41][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane26_strm1_ready         ( DownstreamStackBusLane[41][26].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane26_strm1_cntl          ( DownstreamStackBusLane[41][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane26_strm1_data          ( DownstreamStackBusLane[41][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane26_strm1_data_valid    ( DownstreamStackBusLane[41][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane27_strm0_ready         ( DownstreamStackBusLane[41][27].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane27_strm0_cntl          ( DownstreamStackBusLane[41][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane27_strm0_data          ( DownstreamStackBusLane[41][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane27_strm0_data_valid    ( DownstreamStackBusLane[41][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane27_strm1_ready         ( DownstreamStackBusLane[41][27].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane27_strm1_cntl          ( DownstreamStackBusLane[41][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane27_strm1_data          ( DownstreamStackBusLane[41][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane27_strm1_data_valid    ( DownstreamStackBusLane[41][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane28_strm0_ready         ( DownstreamStackBusLane[41][28].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane28_strm0_cntl          ( DownstreamStackBusLane[41][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane28_strm0_data          ( DownstreamStackBusLane[41][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane28_strm0_data_valid    ( DownstreamStackBusLane[41][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane28_strm1_ready         ( DownstreamStackBusLane[41][28].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane28_strm1_cntl          ( DownstreamStackBusLane[41][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane28_strm1_data          ( DownstreamStackBusLane[41][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane28_strm1_data_valid    ( DownstreamStackBusLane[41][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane29_strm0_ready         ( DownstreamStackBusLane[41][29].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane29_strm0_cntl          ( DownstreamStackBusLane[41][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane29_strm0_data          ( DownstreamStackBusLane[41][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane29_strm0_data_valid    ( DownstreamStackBusLane[41][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane29_strm1_ready         ( DownstreamStackBusLane[41][29].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane29_strm1_cntl          ( DownstreamStackBusLane[41][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane29_strm1_data          ( DownstreamStackBusLane[41][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane29_strm1_data_valid    ( DownstreamStackBusLane[41][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane30_strm0_ready         ( DownstreamStackBusLane[41][30].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane30_strm0_cntl          ( DownstreamStackBusLane[41][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane30_strm0_data          ( DownstreamStackBusLane[41][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane30_strm0_data_valid    ( DownstreamStackBusLane[41][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane30_strm1_ready         ( DownstreamStackBusLane[41][30].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane30_strm1_cntl          ( DownstreamStackBusLane[41][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane30_strm1_data          ( DownstreamStackBusLane[41][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane30_strm1_data_valid    ( DownstreamStackBusLane[41][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 41, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane31_strm0_ready         ( DownstreamStackBusLane[41][31].pe__std__lane_strm0_ready              ),      
        .std__pe41__lane31_strm0_cntl          ( DownstreamStackBusLane[41][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe41__lane31_strm0_data          ( DownstreamStackBusLane[41][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe41__lane31_strm0_data_valid    ( DownstreamStackBusLane[41][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__std__lane31_strm1_ready         ( DownstreamStackBusLane[41][31].pe__std__lane_strm1_ready              ),      
        .std__pe41__lane31_strm1_cntl          ( DownstreamStackBusLane[41][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe41__lane31_strm1_data          ( DownstreamStackBusLane[41][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe41__lane31_strm1_data_valid    ( DownstreamStackBusLane[41][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane0_strm0_ready         ( DownstreamStackBusLane[42][0].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane0_strm0_cntl          ( DownstreamStackBusLane[42][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane0_strm0_data          ( DownstreamStackBusLane[42][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane0_strm0_data_valid    ( DownstreamStackBusLane[42][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane0_strm1_ready         ( DownstreamStackBusLane[42][0].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane0_strm1_cntl          ( DownstreamStackBusLane[42][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane0_strm1_data          ( DownstreamStackBusLane[42][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane0_strm1_data_valid    ( DownstreamStackBusLane[42][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane1_strm0_ready         ( DownstreamStackBusLane[42][1].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane1_strm0_cntl          ( DownstreamStackBusLane[42][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane1_strm0_data          ( DownstreamStackBusLane[42][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane1_strm0_data_valid    ( DownstreamStackBusLane[42][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane1_strm1_ready         ( DownstreamStackBusLane[42][1].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane1_strm1_cntl          ( DownstreamStackBusLane[42][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane1_strm1_data          ( DownstreamStackBusLane[42][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane1_strm1_data_valid    ( DownstreamStackBusLane[42][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane2_strm0_ready         ( DownstreamStackBusLane[42][2].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane2_strm0_cntl          ( DownstreamStackBusLane[42][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane2_strm0_data          ( DownstreamStackBusLane[42][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane2_strm0_data_valid    ( DownstreamStackBusLane[42][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane2_strm1_ready         ( DownstreamStackBusLane[42][2].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane2_strm1_cntl          ( DownstreamStackBusLane[42][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane2_strm1_data          ( DownstreamStackBusLane[42][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane2_strm1_data_valid    ( DownstreamStackBusLane[42][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane3_strm0_ready         ( DownstreamStackBusLane[42][3].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane3_strm0_cntl          ( DownstreamStackBusLane[42][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane3_strm0_data          ( DownstreamStackBusLane[42][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane3_strm0_data_valid    ( DownstreamStackBusLane[42][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane3_strm1_ready         ( DownstreamStackBusLane[42][3].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane3_strm1_cntl          ( DownstreamStackBusLane[42][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane3_strm1_data          ( DownstreamStackBusLane[42][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane3_strm1_data_valid    ( DownstreamStackBusLane[42][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane4_strm0_ready         ( DownstreamStackBusLane[42][4].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane4_strm0_cntl          ( DownstreamStackBusLane[42][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane4_strm0_data          ( DownstreamStackBusLane[42][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane4_strm0_data_valid    ( DownstreamStackBusLane[42][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane4_strm1_ready         ( DownstreamStackBusLane[42][4].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane4_strm1_cntl          ( DownstreamStackBusLane[42][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane4_strm1_data          ( DownstreamStackBusLane[42][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane4_strm1_data_valid    ( DownstreamStackBusLane[42][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane5_strm0_ready         ( DownstreamStackBusLane[42][5].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane5_strm0_cntl          ( DownstreamStackBusLane[42][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane5_strm0_data          ( DownstreamStackBusLane[42][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane5_strm0_data_valid    ( DownstreamStackBusLane[42][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane5_strm1_ready         ( DownstreamStackBusLane[42][5].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane5_strm1_cntl          ( DownstreamStackBusLane[42][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane5_strm1_data          ( DownstreamStackBusLane[42][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane5_strm1_data_valid    ( DownstreamStackBusLane[42][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane6_strm0_ready         ( DownstreamStackBusLane[42][6].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane6_strm0_cntl          ( DownstreamStackBusLane[42][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane6_strm0_data          ( DownstreamStackBusLane[42][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane6_strm0_data_valid    ( DownstreamStackBusLane[42][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane6_strm1_ready         ( DownstreamStackBusLane[42][6].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane6_strm1_cntl          ( DownstreamStackBusLane[42][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane6_strm1_data          ( DownstreamStackBusLane[42][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane6_strm1_data_valid    ( DownstreamStackBusLane[42][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane7_strm0_ready         ( DownstreamStackBusLane[42][7].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane7_strm0_cntl          ( DownstreamStackBusLane[42][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane7_strm0_data          ( DownstreamStackBusLane[42][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane7_strm0_data_valid    ( DownstreamStackBusLane[42][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane7_strm1_ready         ( DownstreamStackBusLane[42][7].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane7_strm1_cntl          ( DownstreamStackBusLane[42][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane7_strm1_data          ( DownstreamStackBusLane[42][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane7_strm1_data_valid    ( DownstreamStackBusLane[42][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane8_strm0_ready         ( DownstreamStackBusLane[42][8].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane8_strm0_cntl          ( DownstreamStackBusLane[42][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane8_strm0_data          ( DownstreamStackBusLane[42][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane8_strm0_data_valid    ( DownstreamStackBusLane[42][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane8_strm1_ready         ( DownstreamStackBusLane[42][8].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane8_strm1_cntl          ( DownstreamStackBusLane[42][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane8_strm1_data          ( DownstreamStackBusLane[42][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane8_strm1_data_valid    ( DownstreamStackBusLane[42][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane9_strm0_ready         ( DownstreamStackBusLane[42][9].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane9_strm0_cntl          ( DownstreamStackBusLane[42][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane9_strm0_data          ( DownstreamStackBusLane[42][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane9_strm0_data_valid    ( DownstreamStackBusLane[42][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane9_strm1_ready         ( DownstreamStackBusLane[42][9].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane9_strm1_cntl          ( DownstreamStackBusLane[42][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane9_strm1_data          ( DownstreamStackBusLane[42][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane9_strm1_data_valid    ( DownstreamStackBusLane[42][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane10_strm0_ready         ( DownstreamStackBusLane[42][10].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane10_strm0_cntl          ( DownstreamStackBusLane[42][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane10_strm0_data          ( DownstreamStackBusLane[42][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane10_strm0_data_valid    ( DownstreamStackBusLane[42][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane10_strm1_ready         ( DownstreamStackBusLane[42][10].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane10_strm1_cntl          ( DownstreamStackBusLane[42][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane10_strm1_data          ( DownstreamStackBusLane[42][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane10_strm1_data_valid    ( DownstreamStackBusLane[42][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane11_strm0_ready         ( DownstreamStackBusLane[42][11].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane11_strm0_cntl          ( DownstreamStackBusLane[42][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane11_strm0_data          ( DownstreamStackBusLane[42][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane11_strm0_data_valid    ( DownstreamStackBusLane[42][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane11_strm1_ready         ( DownstreamStackBusLane[42][11].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane11_strm1_cntl          ( DownstreamStackBusLane[42][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane11_strm1_data          ( DownstreamStackBusLane[42][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane11_strm1_data_valid    ( DownstreamStackBusLane[42][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane12_strm0_ready         ( DownstreamStackBusLane[42][12].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane12_strm0_cntl          ( DownstreamStackBusLane[42][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane12_strm0_data          ( DownstreamStackBusLane[42][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane12_strm0_data_valid    ( DownstreamStackBusLane[42][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane12_strm1_ready         ( DownstreamStackBusLane[42][12].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane12_strm1_cntl          ( DownstreamStackBusLane[42][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane12_strm1_data          ( DownstreamStackBusLane[42][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane12_strm1_data_valid    ( DownstreamStackBusLane[42][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane13_strm0_ready         ( DownstreamStackBusLane[42][13].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane13_strm0_cntl          ( DownstreamStackBusLane[42][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane13_strm0_data          ( DownstreamStackBusLane[42][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane13_strm0_data_valid    ( DownstreamStackBusLane[42][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane13_strm1_ready         ( DownstreamStackBusLane[42][13].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane13_strm1_cntl          ( DownstreamStackBusLane[42][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane13_strm1_data          ( DownstreamStackBusLane[42][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane13_strm1_data_valid    ( DownstreamStackBusLane[42][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane14_strm0_ready         ( DownstreamStackBusLane[42][14].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane14_strm0_cntl          ( DownstreamStackBusLane[42][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane14_strm0_data          ( DownstreamStackBusLane[42][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane14_strm0_data_valid    ( DownstreamStackBusLane[42][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane14_strm1_ready         ( DownstreamStackBusLane[42][14].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane14_strm1_cntl          ( DownstreamStackBusLane[42][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane14_strm1_data          ( DownstreamStackBusLane[42][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane14_strm1_data_valid    ( DownstreamStackBusLane[42][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane15_strm0_ready         ( DownstreamStackBusLane[42][15].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane15_strm0_cntl          ( DownstreamStackBusLane[42][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane15_strm0_data          ( DownstreamStackBusLane[42][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane15_strm0_data_valid    ( DownstreamStackBusLane[42][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane15_strm1_ready         ( DownstreamStackBusLane[42][15].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane15_strm1_cntl          ( DownstreamStackBusLane[42][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane15_strm1_data          ( DownstreamStackBusLane[42][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane15_strm1_data_valid    ( DownstreamStackBusLane[42][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane16_strm0_ready         ( DownstreamStackBusLane[42][16].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane16_strm0_cntl          ( DownstreamStackBusLane[42][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane16_strm0_data          ( DownstreamStackBusLane[42][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane16_strm0_data_valid    ( DownstreamStackBusLane[42][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane16_strm1_ready         ( DownstreamStackBusLane[42][16].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane16_strm1_cntl          ( DownstreamStackBusLane[42][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane16_strm1_data          ( DownstreamStackBusLane[42][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane16_strm1_data_valid    ( DownstreamStackBusLane[42][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane17_strm0_ready         ( DownstreamStackBusLane[42][17].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane17_strm0_cntl          ( DownstreamStackBusLane[42][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane17_strm0_data          ( DownstreamStackBusLane[42][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane17_strm0_data_valid    ( DownstreamStackBusLane[42][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane17_strm1_ready         ( DownstreamStackBusLane[42][17].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane17_strm1_cntl          ( DownstreamStackBusLane[42][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane17_strm1_data          ( DownstreamStackBusLane[42][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane17_strm1_data_valid    ( DownstreamStackBusLane[42][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane18_strm0_ready         ( DownstreamStackBusLane[42][18].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane18_strm0_cntl          ( DownstreamStackBusLane[42][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane18_strm0_data          ( DownstreamStackBusLane[42][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane18_strm0_data_valid    ( DownstreamStackBusLane[42][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane18_strm1_ready         ( DownstreamStackBusLane[42][18].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane18_strm1_cntl          ( DownstreamStackBusLane[42][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane18_strm1_data          ( DownstreamStackBusLane[42][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane18_strm1_data_valid    ( DownstreamStackBusLane[42][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane19_strm0_ready         ( DownstreamStackBusLane[42][19].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane19_strm0_cntl          ( DownstreamStackBusLane[42][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane19_strm0_data          ( DownstreamStackBusLane[42][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane19_strm0_data_valid    ( DownstreamStackBusLane[42][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane19_strm1_ready         ( DownstreamStackBusLane[42][19].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane19_strm1_cntl          ( DownstreamStackBusLane[42][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane19_strm1_data          ( DownstreamStackBusLane[42][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane19_strm1_data_valid    ( DownstreamStackBusLane[42][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane20_strm0_ready         ( DownstreamStackBusLane[42][20].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane20_strm0_cntl          ( DownstreamStackBusLane[42][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane20_strm0_data          ( DownstreamStackBusLane[42][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane20_strm0_data_valid    ( DownstreamStackBusLane[42][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane20_strm1_ready         ( DownstreamStackBusLane[42][20].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane20_strm1_cntl          ( DownstreamStackBusLane[42][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane20_strm1_data          ( DownstreamStackBusLane[42][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane20_strm1_data_valid    ( DownstreamStackBusLane[42][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane21_strm0_ready         ( DownstreamStackBusLane[42][21].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane21_strm0_cntl          ( DownstreamStackBusLane[42][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane21_strm0_data          ( DownstreamStackBusLane[42][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane21_strm0_data_valid    ( DownstreamStackBusLane[42][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane21_strm1_ready         ( DownstreamStackBusLane[42][21].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane21_strm1_cntl          ( DownstreamStackBusLane[42][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane21_strm1_data          ( DownstreamStackBusLane[42][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane21_strm1_data_valid    ( DownstreamStackBusLane[42][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane22_strm0_ready         ( DownstreamStackBusLane[42][22].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane22_strm0_cntl          ( DownstreamStackBusLane[42][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane22_strm0_data          ( DownstreamStackBusLane[42][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane22_strm0_data_valid    ( DownstreamStackBusLane[42][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane22_strm1_ready         ( DownstreamStackBusLane[42][22].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane22_strm1_cntl          ( DownstreamStackBusLane[42][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane22_strm1_data          ( DownstreamStackBusLane[42][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane22_strm1_data_valid    ( DownstreamStackBusLane[42][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane23_strm0_ready         ( DownstreamStackBusLane[42][23].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane23_strm0_cntl          ( DownstreamStackBusLane[42][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane23_strm0_data          ( DownstreamStackBusLane[42][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane23_strm0_data_valid    ( DownstreamStackBusLane[42][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane23_strm1_ready         ( DownstreamStackBusLane[42][23].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane23_strm1_cntl          ( DownstreamStackBusLane[42][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane23_strm1_data          ( DownstreamStackBusLane[42][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane23_strm1_data_valid    ( DownstreamStackBusLane[42][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane24_strm0_ready         ( DownstreamStackBusLane[42][24].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane24_strm0_cntl          ( DownstreamStackBusLane[42][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane24_strm0_data          ( DownstreamStackBusLane[42][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane24_strm0_data_valid    ( DownstreamStackBusLane[42][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane24_strm1_ready         ( DownstreamStackBusLane[42][24].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane24_strm1_cntl          ( DownstreamStackBusLane[42][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane24_strm1_data          ( DownstreamStackBusLane[42][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane24_strm1_data_valid    ( DownstreamStackBusLane[42][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane25_strm0_ready         ( DownstreamStackBusLane[42][25].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane25_strm0_cntl          ( DownstreamStackBusLane[42][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane25_strm0_data          ( DownstreamStackBusLane[42][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane25_strm0_data_valid    ( DownstreamStackBusLane[42][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane25_strm1_ready         ( DownstreamStackBusLane[42][25].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane25_strm1_cntl          ( DownstreamStackBusLane[42][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane25_strm1_data          ( DownstreamStackBusLane[42][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane25_strm1_data_valid    ( DownstreamStackBusLane[42][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane26_strm0_ready         ( DownstreamStackBusLane[42][26].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane26_strm0_cntl          ( DownstreamStackBusLane[42][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane26_strm0_data          ( DownstreamStackBusLane[42][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane26_strm0_data_valid    ( DownstreamStackBusLane[42][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane26_strm1_ready         ( DownstreamStackBusLane[42][26].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane26_strm1_cntl          ( DownstreamStackBusLane[42][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane26_strm1_data          ( DownstreamStackBusLane[42][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane26_strm1_data_valid    ( DownstreamStackBusLane[42][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane27_strm0_ready         ( DownstreamStackBusLane[42][27].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane27_strm0_cntl          ( DownstreamStackBusLane[42][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane27_strm0_data          ( DownstreamStackBusLane[42][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane27_strm0_data_valid    ( DownstreamStackBusLane[42][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane27_strm1_ready         ( DownstreamStackBusLane[42][27].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane27_strm1_cntl          ( DownstreamStackBusLane[42][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane27_strm1_data          ( DownstreamStackBusLane[42][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane27_strm1_data_valid    ( DownstreamStackBusLane[42][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane28_strm0_ready         ( DownstreamStackBusLane[42][28].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane28_strm0_cntl          ( DownstreamStackBusLane[42][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane28_strm0_data          ( DownstreamStackBusLane[42][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane28_strm0_data_valid    ( DownstreamStackBusLane[42][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane28_strm1_ready         ( DownstreamStackBusLane[42][28].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane28_strm1_cntl          ( DownstreamStackBusLane[42][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane28_strm1_data          ( DownstreamStackBusLane[42][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane28_strm1_data_valid    ( DownstreamStackBusLane[42][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane29_strm0_ready         ( DownstreamStackBusLane[42][29].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane29_strm0_cntl          ( DownstreamStackBusLane[42][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane29_strm0_data          ( DownstreamStackBusLane[42][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane29_strm0_data_valid    ( DownstreamStackBusLane[42][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane29_strm1_ready         ( DownstreamStackBusLane[42][29].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane29_strm1_cntl          ( DownstreamStackBusLane[42][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane29_strm1_data          ( DownstreamStackBusLane[42][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane29_strm1_data_valid    ( DownstreamStackBusLane[42][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane30_strm0_ready         ( DownstreamStackBusLane[42][30].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane30_strm0_cntl          ( DownstreamStackBusLane[42][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane30_strm0_data          ( DownstreamStackBusLane[42][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane30_strm0_data_valid    ( DownstreamStackBusLane[42][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane30_strm1_ready         ( DownstreamStackBusLane[42][30].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane30_strm1_cntl          ( DownstreamStackBusLane[42][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane30_strm1_data          ( DownstreamStackBusLane[42][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane30_strm1_data_valid    ( DownstreamStackBusLane[42][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 42, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane31_strm0_ready         ( DownstreamStackBusLane[42][31].pe__std__lane_strm0_ready              ),      
        .std__pe42__lane31_strm0_cntl          ( DownstreamStackBusLane[42][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe42__lane31_strm0_data          ( DownstreamStackBusLane[42][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe42__lane31_strm0_data_valid    ( DownstreamStackBusLane[42][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__std__lane31_strm1_ready         ( DownstreamStackBusLane[42][31].pe__std__lane_strm1_ready              ),      
        .std__pe42__lane31_strm1_cntl          ( DownstreamStackBusLane[42][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe42__lane31_strm1_data          ( DownstreamStackBusLane[42][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe42__lane31_strm1_data_valid    ( DownstreamStackBusLane[42][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane0_strm0_ready         ( DownstreamStackBusLane[43][0].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane0_strm0_cntl          ( DownstreamStackBusLane[43][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane0_strm0_data          ( DownstreamStackBusLane[43][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane0_strm0_data_valid    ( DownstreamStackBusLane[43][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane0_strm1_ready         ( DownstreamStackBusLane[43][0].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane0_strm1_cntl          ( DownstreamStackBusLane[43][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane0_strm1_data          ( DownstreamStackBusLane[43][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane0_strm1_data_valid    ( DownstreamStackBusLane[43][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane1_strm0_ready         ( DownstreamStackBusLane[43][1].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane1_strm0_cntl          ( DownstreamStackBusLane[43][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane1_strm0_data          ( DownstreamStackBusLane[43][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane1_strm0_data_valid    ( DownstreamStackBusLane[43][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane1_strm1_ready         ( DownstreamStackBusLane[43][1].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane1_strm1_cntl          ( DownstreamStackBusLane[43][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane1_strm1_data          ( DownstreamStackBusLane[43][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane1_strm1_data_valid    ( DownstreamStackBusLane[43][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane2_strm0_ready         ( DownstreamStackBusLane[43][2].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane2_strm0_cntl          ( DownstreamStackBusLane[43][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane2_strm0_data          ( DownstreamStackBusLane[43][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane2_strm0_data_valid    ( DownstreamStackBusLane[43][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane2_strm1_ready         ( DownstreamStackBusLane[43][2].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane2_strm1_cntl          ( DownstreamStackBusLane[43][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane2_strm1_data          ( DownstreamStackBusLane[43][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane2_strm1_data_valid    ( DownstreamStackBusLane[43][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane3_strm0_ready         ( DownstreamStackBusLane[43][3].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane3_strm0_cntl          ( DownstreamStackBusLane[43][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane3_strm0_data          ( DownstreamStackBusLane[43][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane3_strm0_data_valid    ( DownstreamStackBusLane[43][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane3_strm1_ready         ( DownstreamStackBusLane[43][3].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane3_strm1_cntl          ( DownstreamStackBusLane[43][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane3_strm1_data          ( DownstreamStackBusLane[43][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane3_strm1_data_valid    ( DownstreamStackBusLane[43][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane4_strm0_ready         ( DownstreamStackBusLane[43][4].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane4_strm0_cntl          ( DownstreamStackBusLane[43][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane4_strm0_data          ( DownstreamStackBusLane[43][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane4_strm0_data_valid    ( DownstreamStackBusLane[43][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane4_strm1_ready         ( DownstreamStackBusLane[43][4].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane4_strm1_cntl          ( DownstreamStackBusLane[43][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane4_strm1_data          ( DownstreamStackBusLane[43][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane4_strm1_data_valid    ( DownstreamStackBusLane[43][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane5_strm0_ready         ( DownstreamStackBusLane[43][5].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane5_strm0_cntl          ( DownstreamStackBusLane[43][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane5_strm0_data          ( DownstreamStackBusLane[43][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane5_strm0_data_valid    ( DownstreamStackBusLane[43][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane5_strm1_ready         ( DownstreamStackBusLane[43][5].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane5_strm1_cntl          ( DownstreamStackBusLane[43][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane5_strm1_data          ( DownstreamStackBusLane[43][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane5_strm1_data_valid    ( DownstreamStackBusLane[43][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane6_strm0_ready         ( DownstreamStackBusLane[43][6].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane6_strm0_cntl          ( DownstreamStackBusLane[43][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane6_strm0_data          ( DownstreamStackBusLane[43][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane6_strm0_data_valid    ( DownstreamStackBusLane[43][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane6_strm1_ready         ( DownstreamStackBusLane[43][6].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane6_strm1_cntl          ( DownstreamStackBusLane[43][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane6_strm1_data          ( DownstreamStackBusLane[43][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane6_strm1_data_valid    ( DownstreamStackBusLane[43][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane7_strm0_ready         ( DownstreamStackBusLane[43][7].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane7_strm0_cntl          ( DownstreamStackBusLane[43][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane7_strm0_data          ( DownstreamStackBusLane[43][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane7_strm0_data_valid    ( DownstreamStackBusLane[43][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane7_strm1_ready         ( DownstreamStackBusLane[43][7].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane7_strm1_cntl          ( DownstreamStackBusLane[43][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane7_strm1_data          ( DownstreamStackBusLane[43][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane7_strm1_data_valid    ( DownstreamStackBusLane[43][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane8_strm0_ready         ( DownstreamStackBusLane[43][8].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane8_strm0_cntl          ( DownstreamStackBusLane[43][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane8_strm0_data          ( DownstreamStackBusLane[43][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane8_strm0_data_valid    ( DownstreamStackBusLane[43][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane8_strm1_ready         ( DownstreamStackBusLane[43][8].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane8_strm1_cntl          ( DownstreamStackBusLane[43][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane8_strm1_data          ( DownstreamStackBusLane[43][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane8_strm1_data_valid    ( DownstreamStackBusLane[43][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane9_strm0_ready         ( DownstreamStackBusLane[43][9].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane9_strm0_cntl          ( DownstreamStackBusLane[43][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane9_strm0_data          ( DownstreamStackBusLane[43][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane9_strm0_data_valid    ( DownstreamStackBusLane[43][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane9_strm1_ready         ( DownstreamStackBusLane[43][9].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane9_strm1_cntl          ( DownstreamStackBusLane[43][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane9_strm1_data          ( DownstreamStackBusLane[43][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane9_strm1_data_valid    ( DownstreamStackBusLane[43][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane10_strm0_ready         ( DownstreamStackBusLane[43][10].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane10_strm0_cntl          ( DownstreamStackBusLane[43][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane10_strm0_data          ( DownstreamStackBusLane[43][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane10_strm0_data_valid    ( DownstreamStackBusLane[43][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane10_strm1_ready         ( DownstreamStackBusLane[43][10].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane10_strm1_cntl          ( DownstreamStackBusLane[43][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane10_strm1_data          ( DownstreamStackBusLane[43][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane10_strm1_data_valid    ( DownstreamStackBusLane[43][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane11_strm0_ready         ( DownstreamStackBusLane[43][11].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane11_strm0_cntl          ( DownstreamStackBusLane[43][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane11_strm0_data          ( DownstreamStackBusLane[43][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane11_strm0_data_valid    ( DownstreamStackBusLane[43][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane11_strm1_ready         ( DownstreamStackBusLane[43][11].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane11_strm1_cntl          ( DownstreamStackBusLane[43][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane11_strm1_data          ( DownstreamStackBusLane[43][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane11_strm1_data_valid    ( DownstreamStackBusLane[43][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane12_strm0_ready         ( DownstreamStackBusLane[43][12].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane12_strm0_cntl          ( DownstreamStackBusLane[43][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane12_strm0_data          ( DownstreamStackBusLane[43][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane12_strm0_data_valid    ( DownstreamStackBusLane[43][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane12_strm1_ready         ( DownstreamStackBusLane[43][12].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane12_strm1_cntl          ( DownstreamStackBusLane[43][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane12_strm1_data          ( DownstreamStackBusLane[43][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane12_strm1_data_valid    ( DownstreamStackBusLane[43][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane13_strm0_ready         ( DownstreamStackBusLane[43][13].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane13_strm0_cntl          ( DownstreamStackBusLane[43][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane13_strm0_data          ( DownstreamStackBusLane[43][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane13_strm0_data_valid    ( DownstreamStackBusLane[43][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane13_strm1_ready         ( DownstreamStackBusLane[43][13].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane13_strm1_cntl          ( DownstreamStackBusLane[43][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane13_strm1_data          ( DownstreamStackBusLane[43][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane13_strm1_data_valid    ( DownstreamStackBusLane[43][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane14_strm0_ready         ( DownstreamStackBusLane[43][14].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane14_strm0_cntl          ( DownstreamStackBusLane[43][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane14_strm0_data          ( DownstreamStackBusLane[43][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane14_strm0_data_valid    ( DownstreamStackBusLane[43][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane14_strm1_ready         ( DownstreamStackBusLane[43][14].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane14_strm1_cntl          ( DownstreamStackBusLane[43][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane14_strm1_data          ( DownstreamStackBusLane[43][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane14_strm1_data_valid    ( DownstreamStackBusLane[43][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane15_strm0_ready         ( DownstreamStackBusLane[43][15].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane15_strm0_cntl          ( DownstreamStackBusLane[43][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane15_strm0_data          ( DownstreamStackBusLane[43][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane15_strm0_data_valid    ( DownstreamStackBusLane[43][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane15_strm1_ready         ( DownstreamStackBusLane[43][15].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane15_strm1_cntl          ( DownstreamStackBusLane[43][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane15_strm1_data          ( DownstreamStackBusLane[43][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane15_strm1_data_valid    ( DownstreamStackBusLane[43][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane16_strm0_ready         ( DownstreamStackBusLane[43][16].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane16_strm0_cntl          ( DownstreamStackBusLane[43][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane16_strm0_data          ( DownstreamStackBusLane[43][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane16_strm0_data_valid    ( DownstreamStackBusLane[43][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane16_strm1_ready         ( DownstreamStackBusLane[43][16].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane16_strm1_cntl          ( DownstreamStackBusLane[43][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane16_strm1_data          ( DownstreamStackBusLane[43][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane16_strm1_data_valid    ( DownstreamStackBusLane[43][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane17_strm0_ready         ( DownstreamStackBusLane[43][17].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane17_strm0_cntl          ( DownstreamStackBusLane[43][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane17_strm0_data          ( DownstreamStackBusLane[43][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane17_strm0_data_valid    ( DownstreamStackBusLane[43][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane17_strm1_ready         ( DownstreamStackBusLane[43][17].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane17_strm1_cntl          ( DownstreamStackBusLane[43][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane17_strm1_data          ( DownstreamStackBusLane[43][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane17_strm1_data_valid    ( DownstreamStackBusLane[43][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane18_strm0_ready         ( DownstreamStackBusLane[43][18].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane18_strm0_cntl          ( DownstreamStackBusLane[43][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane18_strm0_data          ( DownstreamStackBusLane[43][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane18_strm0_data_valid    ( DownstreamStackBusLane[43][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane18_strm1_ready         ( DownstreamStackBusLane[43][18].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane18_strm1_cntl          ( DownstreamStackBusLane[43][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane18_strm1_data          ( DownstreamStackBusLane[43][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane18_strm1_data_valid    ( DownstreamStackBusLane[43][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane19_strm0_ready         ( DownstreamStackBusLane[43][19].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane19_strm0_cntl          ( DownstreamStackBusLane[43][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane19_strm0_data          ( DownstreamStackBusLane[43][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane19_strm0_data_valid    ( DownstreamStackBusLane[43][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane19_strm1_ready         ( DownstreamStackBusLane[43][19].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane19_strm1_cntl          ( DownstreamStackBusLane[43][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane19_strm1_data          ( DownstreamStackBusLane[43][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane19_strm1_data_valid    ( DownstreamStackBusLane[43][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane20_strm0_ready         ( DownstreamStackBusLane[43][20].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane20_strm0_cntl          ( DownstreamStackBusLane[43][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane20_strm0_data          ( DownstreamStackBusLane[43][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane20_strm0_data_valid    ( DownstreamStackBusLane[43][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane20_strm1_ready         ( DownstreamStackBusLane[43][20].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane20_strm1_cntl          ( DownstreamStackBusLane[43][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane20_strm1_data          ( DownstreamStackBusLane[43][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane20_strm1_data_valid    ( DownstreamStackBusLane[43][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane21_strm0_ready         ( DownstreamStackBusLane[43][21].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane21_strm0_cntl          ( DownstreamStackBusLane[43][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane21_strm0_data          ( DownstreamStackBusLane[43][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane21_strm0_data_valid    ( DownstreamStackBusLane[43][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane21_strm1_ready         ( DownstreamStackBusLane[43][21].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane21_strm1_cntl          ( DownstreamStackBusLane[43][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane21_strm1_data          ( DownstreamStackBusLane[43][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane21_strm1_data_valid    ( DownstreamStackBusLane[43][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane22_strm0_ready         ( DownstreamStackBusLane[43][22].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane22_strm0_cntl          ( DownstreamStackBusLane[43][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane22_strm0_data          ( DownstreamStackBusLane[43][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane22_strm0_data_valid    ( DownstreamStackBusLane[43][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane22_strm1_ready         ( DownstreamStackBusLane[43][22].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane22_strm1_cntl          ( DownstreamStackBusLane[43][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane22_strm1_data          ( DownstreamStackBusLane[43][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane22_strm1_data_valid    ( DownstreamStackBusLane[43][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane23_strm0_ready         ( DownstreamStackBusLane[43][23].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane23_strm0_cntl          ( DownstreamStackBusLane[43][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane23_strm0_data          ( DownstreamStackBusLane[43][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane23_strm0_data_valid    ( DownstreamStackBusLane[43][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane23_strm1_ready         ( DownstreamStackBusLane[43][23].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane23_strm1_cntl          ( DownstreamStackBusLane[43][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane23_strm1_data          ( DownstreamStackBusLane[43][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane23_strm1_data_valid    ( DownstreamStackBusLane[43][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane24_strm0_ready         ( DownstreamStackBusLane[43][24].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane24_strm0_cntl          ( DownstreamStackBusLane[43][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane24_strm0_data          ( DownstreamStackBusLane[43][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane24_strm0_data_valid    ( DownstreamStackBusLane[43][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane24_strm1_ready         ( DownstreamStackBusLane[43][24].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane24_strm1_cntl          ( DownstreamStackBusLane[43][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane24_strm1_data          ( DownstreamStackBusLane[43][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane24_strm1_data_valid    ( DownstreamStackBusLane[43][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane25_strm0_ready         ( DownstreamStackBusLane[43][25].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane25_strm0_cntl          ( DownstreamStackBusLane[43][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane25_strm0_data          ( DownstreamStackBusLane[43][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane25_strm0_data_valid    ( DownstreamStackBusLane[43][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane25_strm1_ready         ( DownstreamStackBusLane[43][25].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane25_strm1_cntl          ( DownstreamStackBusLane[43][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane25_strm1_data          ( DownstreamStackBusLane[43][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane25_strm1_data_valid    ( DownstreamStackBusLane[43][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane26_strm0_ready         ( DownstreamStackBusLane[43][26].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane26_strm0_cntl          ( DownstreamStackBusLane[43][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane26_strm0_data          ( DownstreamStackBusLane[43][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane26_strm0_data_valid    ( DownstreamStackBusLane[43][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane26_strm1_ready         ( DownstreamStackBusLane[43][26].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane26_strm1_cntl          ( DownstreamStackBusLane[43][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane26_strm1_data          ( DownstreamStackBusLane[43][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane26_strm1_data_valid    ( DownstreamStackBusLane[43][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane27_strm0_ready         ( DownstreamStackBusLane[43][27].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane27_strm0_cntl          ( DownstreamStackBusLane[43][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane27_strm0_data          ( DownstreamStackBusLane[43][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane27_strm0_data_valid    ( DownstreamStackBusLane[43][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane27_strm1_ready         ( DownstreamStackBusLane[43][27].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane27_strm1_cntl          ( DownstreamStackBusLane[43][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane27_strm1_data          ( DownstreamStackBusLane[43][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane27_strm1_data_valid    ( DownstreamStackBusLane[43][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane28_strm0_ready         ( DownstreamStackBusLane[43][28].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane28_strm0_cntl          ( DownstreamStackBusLane[43][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane28_strm0_data          ( DownstreamStackBusLane[43][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane28_strm0_data_valid    ( DownstreamStackBusLane[43][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane28_strm1_ready         ( DownstreamStackBusLane[43][28].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane28_strm1_cntl          ( DownstreamStackBusLane[43][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane28_strm1_data          ( DownstreamStackBusLane[43][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane28_strm1_data_valid    ( DownstreamStackBusLane[43][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane29_strm0_ready         ( DownstreamStackBusLane[43][29].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane29_strm0_cntl          ( DownstreamStackBusLane[43][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane29_strm0_data          ( DownstreamStackBusLane[43][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane29_strm0_data_valid    ( DownstreamStackBusLane[43][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane29_strm1_ready         ( DownstreamStackBusLane[43][29].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane29_strm1_cntl          ( DownstreamStackBusLane[43][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane29_strm1_data          ( DownstreamStackBusLane[43][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane29_strm1_data_valid    ( DownstreamStackBusLane[43][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane30_strm0_ready         ( DownstreamStackBusLane[43][30].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane30_strm0_cntl          ( DownstreamStackBusLane[43][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane30_strm0_data          ( DownstreamStackBusLane[43][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane30_strm0_data_valid    ( DownstreamStackBusLane[43][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane30_strm1_ready         ( DownstreamStackBusLane[43][30].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane30_strm1_cntl          ( DownstreamStackBusLane[43][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane30_strm1_data          ( DownstreamStackBusLane[43][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane30_strm1_data_valid    ( DownstreamStackBusLane[43][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 43, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane31_strm0_ready         ( DownstreamStackBusLane[43][31].pe__std__lane_strm0_ready              ),      
        .std__pe43__lane31_strm0_cntl          ( DownstreamStackBusLane[43][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe43__lane31_strm0_data          ( DownstreamStackBusLane[43][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe43__lane31_strm0_data_valid    ( DownstreamStackBusLane[43][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__std__lane31_strm1_ready         ( DownstreamStackBusLane[43][31].pe__std__lane_strm1_ready              ),      
        .std__pe43__lane31_strm1_cntl          ( DownstreamStackBusLane[43][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe43__lane31_strm1_data          ( DownstreamStackBusLane[43][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe43__lane31_strm1_data_valid    ( DownstreamStackBusLane[43][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane0_strm0_ready         ( DownstreamStackBusLane[44][0].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane0_strm0_cntl          ( DownstreamStackBusLane[44][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane0_strm0_data          ( DownstreamStackBusLane[44][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane0_strm0_data_valid    ( DownstreamStackBusLane[44][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane0_strm1_ready         ( DownstreamStackBusLane[44][0].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane0_strm1_cntl          ( DownstreamStackBusLane[44][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane0_strm1_data          ( DownstreamStackBusLane[44][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane0_strm1_data_valid    ( DownstreamStackBusLane[44][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane1_strm0_ready         ( DownstreamStackBusLane[44][1].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane1_strm0_cntl          ( DownstreamStackBusLane[44][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane1_strm0_data          ( DownstreamStackBusLane[44][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane1_strm0_data_valid    ( DownstreamStackBusLane[44][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane1_strm1_ready         ( DownstreamStackBusLane[44][1].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane1_strm1_cntl          ( DownstreamStackBusLane[44][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane1_strm1_data          ( DownstreamStackBusLane[44][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane1_strm1_data_valid    ( DownstreamStackBusLane[44][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane2_strm0_ready         ( DownstreamStackBusLane[44][2].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane2_strm0_cntl          ( DownstreamStackBusLane[44][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane2_strm0_data          ( DownstreamStackBusLane[44][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane2_strm0_data_valid    ( DownstreamStackBusLane[44][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane2_strm1_ready         ( DownstreamStackBusLane[44][2].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane2_strm1_cntl          ( DownstreamStackBusLane[44][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane2_strm1_data          ( DownstreamStackBusLane[44][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane2_strm1_data_valid    ( DownstreamStackBusLane[44][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane3_strm0_ready         ( DownstreamStackBusLane[44][3].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane3_strm0_cntl          ( DownstreamStackBusLane[44][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane3_strm0_data          ( DownstreamStackBusLane[44][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane3_strm0_data_valid    ( DownstreamStackBusLane[44][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane3_strm1_ready         ( DownstreamStackBusLane[44][3].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane3_strm1_cntl          ( DownstreamStackBusLane[44][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane3_strm1_data          ( DownstreamStackBusLane[44][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane3_strm1_data_valid    ( DownstreamStackBusLane[44][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane4_strm0_ready         ( DownstreamStackBusLane[44][4].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane4_strm0_cntl          ( DownstreamStackBusLane[44][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane4_strm0_data          ( DownstreamStackBusLane[44][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane4_strm0_data_valid    ( DownstreamStackBusLane[44][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane4_strm1_ready         ( DownstreamStackBusLane[44][4].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane4_strm1_cntl          ( DownstreamStackBusLane[44][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane4_strm1_data          ( DownstreamStackBusLane[44][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane4_strm1_data_valid    ( DownstreamStackBusLane[44][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane5_strm0_ready         ( DownstreamStackBusLane[44][5].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane5_strm0_cntl          ( DownstreamStackBusLane[44][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane5_strm0_data          ( DownstreamStackBusLane[44][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane5_strm0_data_valid    ( DownstreamStackBusLane[44][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane5_strm1_ready         ( DownstreamStackBusLane[44][5].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane5_strm1_cntl          ( DownstreamStackBusLane[44][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane5_strm1_data          ( DownstreamStackBusLane[44][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane5_strm1_data_valid    ( DownstreamStackBusLane[44][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane6_strm0_ready         ( DownstreamStackBusLane[44][6].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane6_strm0_cntl          ( DownstreamStackBusLane[44][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane6_strm0_data          ( DownstreamStackBusLane[44][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane6_strm0_data_valid    ( DownstreamStackBusLane[44][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane6_strm1_ready         ( DownstreamStackBusLane[44][6].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane6_strm1_cntl          ( DownstreamStackBusLane[44][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane6_strm1_data          ( DownstreamStackBusLane[44][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane6_strm1_data_valid    ( DownstreamStackBusLane[44][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane7_strm0_ready         ( DownstreamStackBusLane[44][7].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane7_strm0_cntl          ( DownstreamStackBusLane[44][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane7_strm0_data          ( DownstreamStackBusLane[44][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane7_strm0_data_valid    ( DownstreamStackBusLane[44][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane7_strm1_ready         ( DownstreamStackBusLane[44][7].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane7_strm1_cntl          ( DownstreamStackBusLane[44][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane7_strm1_data          ( DownstreamStackBusLane[44][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane7_strm1_data_valid    ( DownstreamStackBusLane[44][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane8_strm0_ready         ( DownstreamStackBusLane[44][8].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane8_strm0_cntl          ( DownstreamStackBusLane[44][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane8_strm0_data          ( DownstreamStackBusLane[44][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane8_strm0_data_valid    ( DownstreamStackBusLane[44][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane8_strm1_ready         ( DownstreamStackBusLane[44][8].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane8_strm1_cntl          ( DownstreamStackBusLane[44][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane8_strm1_data          ( DownstreamStackBusLane[44][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane8_strm1_data_valid    ( DownstreamStackBusLane[44][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane9_strm0_ready         ( DownstreamStackBusLane[44][9].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane9_strm0_cntl          ( DownstreamStackBusLane[44][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane9_strm0_data          ( DownstreamStackBusLane[44][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane9_strm0_data_valid    ( DownstreamStackBusLane[44][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane9_strm1_ready         ( DownstreamStackBusLane[44][9].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane9_strm1_cntl          ( DownstreamStackBusLane[44][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane9_strm1_data          ( DownstreamStackBusLane[44][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane9_strm1_data_valid    ( DownstreamStackBusLane[44][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane10_strm0_ready         ( DownstreamStackBusLane[44][10].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane10_strm0_cntl          ( DownstreamStackBusLane[44][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane10_strm0_data          ( DownstreamStackBusLane[44][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane10_strm0_data_valid    ( DownstreamStackBusLane[44][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane10_strm1_ready         ( DownstreamStackBusLane[44][10].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane10_strm1_cntl          ( DownstreamStackBusLane[44][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane10_strm1_data          ( DownstreamStackBusLane[44][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane10_strm1_data_valid    ( DownstreamStackBusLane[44][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane11_strm0_ready         ( DownstreamStackBusLane[44][11].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane11_strm0_cntl          ( DownstreamStackBusLane[44][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane11_strm0_data          ( DownstreamStackBusLane[44][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane11_strm0_data_valid    ( DownstreamStackBusLane[44][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane11_strm1_ready         ( DownstreamStackBusLane[44][11].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane11_strm1_cntl          ( DownstreamStackBusLane[44][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane11_strm1_data          ( DownstreamStackBusLane[44][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane11_strm1_data_valid    ( DownstreamStackBusLane[44][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane12_strm0_ready         ( DownstreamStackBusLane[44][12].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane12_strm0_cntl          ( DownstreamStackBusLane[44][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane12_strm0_data          ( DownstreamStackBusLane[44][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane12_strm0_data_valid    ( DownstreamStackBusLane[44][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane12_strm1_ready         ( DownstreamStackBusLane[44][12].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane12_strm1_cntl          ( DownstreamStackBusLane[44][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane12_strm1_data          ( DownstreamStackBusLane[44][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane12_strm1_data_valid    ( DownstreamStackBusLane[44][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane13_strm0_ready         ( DownstreamStackBusLane[44][13].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane13_strm0_cntl          ( DownstreamStackBusLane[44][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane13_strm0_data          ( DownstreamStackBusLane[44][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane13_strm0_data_valid    ( DownstreamStackBusLane[44][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane13_strm1_ready         ( DownstreamStackBusLane[44][13].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane13_strm1_cntl          ( DownstreamStackBusLane[44][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane13_strm1_data          ( DownstreamStackBusLane[44][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane13_strm1_data_valid    ( DownstreamStackBusLane[44][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane14_strm0_ready         ( DownstreamStackBusLane[44][14].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane14_strm0_cntl          ( DownstreamStackBusLane[44][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane14_strm0_data          ( DownstreamStackBusLane[44][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane14_strm0_data_valid    ( DownstreamStackBusLane[44][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane14_strm1_ready         ( DownstreamStackBusLane[44][14].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane14_strm1_cntl          ( DownstreamStackBusLane[44][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane14_strm1_data          ( DownstreamStackBusLane[44][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane14_strm1_data_valid    ( DownstreamStackBusLane[44][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane15_strm0_ready         ( DownstreamStackBusLane[44][15].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane15_strm0_cntl          ( DownstreamStackBusLane[44][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane15_strm0_data          ( DownstreamStackBusLane[44][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane15_strm0_data_valid    ( DownstreamStackBusLane[44][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane15_strm1_ready         ( DownstreamStackBusLane[44][15].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane15_strm1_cntl          ( DownstreamStackBusLane[44][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane15_strm1_data          ( DownstreamStackBusLane[44][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane15_strm1_data_valid    ( DownstreamStackBusLane[44][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane16_strm0_ready         ( DownstreamStackBusLane[44][16].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane16_strm0_cntl          ( DownstreamStackBusLane[44][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane16_strm0_data          ( DownstreamStackBusLane[44][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane16_strm0_data_valid    ( DownstreamStackBusLane[44][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane16_strm1_ready         ( DownstreamStackBusLane[44][16].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane16_strm1_cntl          ( DownstreamStackBusLane[44][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane16_strm1_data          ( DownstreamStackBusLane[44][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane16_strm1_data_valid    ( DownstreamStackBusLane[44][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane17_strm0_ready         ( DownstreamStackBusLane[44][17].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane17_strm0_cntl          ( DownstreamStackBusLane[44][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane17_strm0_data          ( DownstreamStackBusLane[44][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane17_strm0_data_valid    ( DownstreamStackBusLane[44][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane17_strm1_ready         ( DownstreamStackBusLane[44][17].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane17_strm1_cntl          ( DownstreamStackBusLane[44][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane17_strm1_data          ( DownstreamStackBusLane[44][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane17_strm1_data_valid    ( DownstreamStackBusLane[44][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane18_strm0_ready         ( DownstreamStackBusLane[44][18].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane18_strm0_cntl          ( DownstreamStackBusLane[44][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane18_strm0_data          ( DownstreamStackBusLane[44][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane18_strm0_data_valid    ( DownstreamStackBusLane[44][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane18_strm1_ready         ( DownstreamStackBusLane[44][18].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane18_strm1_cntl          ( DownstreamStackBusLane[44][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane18_strm1_data          ( DownstreamStackBusLane[44][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane18_strm1_data_valid    ( DownstreamStackBusLane[44][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane19_strm0_ready         ( DownstreamStackBusLane[44][19].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane19_strm0_cntl          ( DownstreamStackBusLane[44][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane19_strm0_data          ( DownstreamStackBusLane[44][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane19_strm0_data_valid    ( DownstreamStackBusLane[44][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane19_strm1_ready         ( DownstreamStackBusLane[44][19].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane19_strm1_cntl          ( DownstreamStackBusLane[44][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane19_strm1_data          ( DownstreamStackBusLane[44][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane19_strm1_data_valid    ( DownstreamStackBusLane[44][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane20_strm0_ready         ( DownstreamStackBusLane[44][20].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane20_strm0_cntl          ( DownstreamStackBusLane[44][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane20_strm0_data          ( DownstreamStackBusLane[44][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane20_strm0_data_valid    ( DownstreamStackBusLane[44][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane20_strm1_ready         ( DownstreamStackBusLane[44][20].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane20_strm1_cntl          ( DownstreamStackBusLane[44][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane20_strm1_data          ( DownstreamStackBusLane[44][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane20_strm1_data_valid    ( DownstreamStackBusLane[44][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane21_strm0_ready         ( DownstreamStackBusLane[44][21].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane21_strm0_cntl          ( DownstreamStackBusLane[44][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane21_strm0_data          ( DownstreamStackBusLane[44][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane21_strm0_data_valid    ( DownstreamStackBusLane[44][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane21_strm1_ready         ( DownstreamStackBusLane[44][21].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane21_strm1_cntl          ( DownstreamStackBusLane[44][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane21_strm1_data          ( DownstreamStackBusLane[44][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane21_strm1_data_valid    ( DownstreamStackBusLane[44][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane22_strm0_ready         ( DownstreamStackBusLane[44][22].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane22_strm0_cntl          ( DownstreamStackBusLane[44][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane22_strm0_data          ( DownstreamStackBusLane[44][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane22_strm0_data_valid    ( DownstreamStackBusLane[44][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane22_strm1_ready         ( DownstreamStackBusLane[44][22].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane22_strm1_cntl          ( DownstreamStackBusLane[44][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane22_strm1_data          ( DownstreamStackBusLane[44][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane22_strm1_data_valid    ( DownstreamStackBusLane[44][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane23_strm0_ready         ( DownstreamStackBusLane[44][23].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane23_strm0_cntl          ( DownstreamStackBusLane[44][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane23_strm0_data          ( DownstreamStackBusLane[44][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane23_strm0_data_valid    ( DownstreamStackBusLane[44][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane23_strm1_ready         ( DownstreamStackBusLane[44][23].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane23_strm1_cntl          ( DownstreamStackBusLane[44][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane23_strm1_data          ( DownstreamStackBusLane[44][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane23_strm1_data_valid    ( DownstreamStackBusLane[44][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane24_strm0_ready         ( DownstreamStackBusLane[44][24].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane24_strm0_cntl          ( DownstreamStackBusLane[44][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane24_strm0_data          ( DownstreamStackBusLane[44][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane24_strm0_data_valid    ( DownstreamStackBusLane[44][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane24_strm1_ready         ( DownstreamStackBusLane[44][24].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane24_strm1_cntl          ( DownstreamStackBusLane[44][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane24_strm1_data          ( DownstreamStackBusLane[44][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane24_strm1_data_valid    ( DownstreamStackBusLane[44][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane25_strm0_ready         ( DownstreamStackBusLane[44][25].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane25_strm0_cntl          ( DownstreamStackBusLane[44][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane25_strm0_data          ( DownstreamStackBusLane[44][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane25_strm0_data_valid    ( DownstreamStackBusLane[44][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane25_strm1_ready         ( DownstreamStackBusLane[44][25].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane25_strm1_cntl          ( DownstreamStackBusLane[44][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane25_strm1_data          ( DownstreamStackBusLane[44][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane25_strm1_data_valid    ( DownstreamStackBusLane[44][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane26_strm0_ready         ( DownstreamStackBusLane[44][26].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane26_strm0_cntl          ( DownstreamStackBusLane[44][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane26_strm0_data          ( DownstreamStackBusLane[44][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane26_strm0_data_valid    ( DownstreamStackBusLane[44][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane26_strm1_ready         ( DownstreamStackBusLane[44][26].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane26_strm1_cntl          ( DownstreamStackBusLane[44][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane26_strm1_data          ( DownstreamStackBusLane[44][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane26_strm1_data_valid    ( DownstreamStackBusLane[44][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane27_strm0_ready         ( DownstreamStackBusLane[44][27].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane27_strm0_cntl          ( DownstreamStackBusLane[44][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane27_strm0_data          ( DownstreamStackBusLane[44][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane27_strm0_data_valid    ( DownstreamStackBusLane[44][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane27_strm1_ready         ( DownstreamStackBusLane[44][27].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane27_strm1_cntl          ( DownstreamStackBusLane[44][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane27_strm1_data          ( DownstreamStackBusLane[44][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane27_strm1_data_valid    ( DownstreamStackBusLane[44][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane28_strm0_ready         ( DownstreamStackBusLane[44][28].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane28_strm0_cntl          ( DownstreamStackBusLane[44][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane28_strm0_data          ( DownstreamStackBusLane[44][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane28_strm0_data_valid    ( DownstreamStackBusLane[44][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane28_strm1_ready         ( DownstreamStackBusLane[44][28].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane28_strm1_cntl          ( DownstreamStackBusLane[44][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane28_strm1_data          ( DownstreamStackBusLane[44][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane28_strm1_data_valid    ( DownstreamStackBusLane[44][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane29_strm0_ready         ( DownstreamStackBusLane[44][29].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane29_strm0_cntl          ( DownstreamStackBusLane[44][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane29_strm0_data          ( DownstreamStackBusLane[44][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane29_strm0_data_valid    ( DownstreamStackBusLane[44][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane29_strm1_ready         ( DownstreamStackBusLane[44][29].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane29_strm1_cntl          ( DownstreamStackBusLane[44][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane29_strm1_data          ( DownstreamStackBusLane[44][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane29_strm1_data_valid    ( DownstreamStackBusLane[44][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane30_strm0_ready         ( DownstreamStackBusLane[44][30].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane30_strm0_cntl          ( DownstreamStackBusLane[44][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane30_strm0_data          ( DownstreamStackBusLane[44][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane30_strm0_data_valid    ( DownstreamStackBusLane[44][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane30_strm1_ready         ( DownstreamStackBusLane[44][30].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane30_strm1_cntl          ( DownstreamStackBusLane[44][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane30_strm1_data          ( DownstreamStackBusLane[44][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane30_strm1_data_valid    ( DownstreamStackBusLane[44][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 44, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane31_strm0_ready         ( DownstreamStackBusLane[44][31].pe__std__lane_strm0_ready              ),      
        .std__pe44__lane31_strm0_cntl          ( DownstreamStackBusLane[44][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe44__lane31_strm0_data          ( DownstreamStackBusLane[44][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe44__lane31_strm0_data_valid    ( DownstreamStackBusLane[44][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__std__lane31_strm1_ready         ( DownstreamStackBusLane[44][31].pe__std__lane_strm1_ready              ),      
        .std__pe44__lane31_strm1_cntl          ( DownstreamStackBusLane[44][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe44__lane31_strm1_data          ( DownstreamStackBusLane[44][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe44__lane31_strm1_data_valid    ( DownstreamStackBusLane[44][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane0_strm0_ready         ( DownstreamStackBusLane[45][0].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane0_strm0_cntl          ( DownstreamStackBusLane[45][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane0_strm0_data          ( DownstreamStackBusLane[45][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane0_strm0_data_valid    ( DownstreamStackBusLane[45][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane0_strm1_ready         ( DownstreamStackBusLane[45][0].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane0_strm1_cntl          ( DownstreamStackBusLane[45][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane0_strm1_data          ( DownstreamStackBusLane[45][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane0_strm1_data_valid    ( DownstreamStackBusLane[45][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane1_strm0_ready         ( DownstreamStackBusLane[45][1].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane1_strm0_cntl          ( DownstreamStackBusLane[45][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane1_strm0_data          ( DownstreamStackBusLane[45][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane1_strm0_data_valid    ( DownstreamStackBusLane[45][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane1_strm1_ready         ( DownstreamStackBusLane[45][1].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane1_strm1_cntl          ( DownstreamStackBusLane[45][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane1_strm1_data          ( DownstreamStackBusLane[45][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane1_strm1_data_valid    ( DownstreamStackBusLane[45][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane2_strm0_ready         ( DownstreamStackBusLane[45][2].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane2_strm0_cntl          ( DownstreamStackBusLane[45][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane2_strm0_data          ( DownstreamStackBusLane[45][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane2_strm0_data_valid    ( DownstreamStackBusLane[45][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane2_strm1_ready         ( DownstreamStackBusLane[45][2].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane2_strm1_cntl          ( DownstreamStackBusLane[45][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane2_strm1_data          ( DownstreamStackBusLane[45][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane2_strm1_data_valid    ( DownstreamStackBusLane[45][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane3_strm0_ready         ( DownstreamStackBusLane[45][3].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane3_strm0_cntl          ( DownstreamStackBusLane[45][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane3_strm0_data          ( DownstreamStackBusLane[45][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane3_strm0_data_valid    ( DownstreamStackBusLane[45][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane3_strm1_ready         ( DownstreamStackBusLane[45][3].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane3_strm1_cntl          ( DownstreamStackBusLane[45][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane3_strm1_data          ( DownstreamStackBusLane[45][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane3_strm1_data_valid    ( DownstreamStackBusLane[45][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane4_strm0_ready         ( DownstreamStackBusLane[45][4].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane4_strm0_cntl          ( DownstreamStackBusLane[45][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane4_strm0_data          ( DownstreamStackBusLane[45][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane4_strm0_data_valid    ( DownstreamStackBusLane[45][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane4_strm1_ready         ( DownstreamStackBusLane[45][4].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane4_strm1_cntl          ( DownstreamStackBusLane[45][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane4_strm1_data          ( DownstreamStackBusLane[45][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane4_strm1_data_valid    ( DownstreamStackBusLane[45][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane5_strm0_ready         ( DownstreamStackBusLane[45][5].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane5_strm0_cntl          ( DownstreamStackBusLane[45][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane5_strm0_data          ( DownstreamStackBusLane[45][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane5_strm0_data_valid    ( DownstreamStackBusLane[45][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane5_strm1_ready         ( DownstreamStackBusLane[45][5].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane5_strm1_cntl          ( DownstreamStackBusLane[45][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane5_strm1_data          ( DownstreamStackBusLane[45][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane5_strm1_data_valid    ( DownstreamStackBusLane[45][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane6_strm0_ready         ( DownstreamStackBusLane[45][6].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane6_strm0_cntl          ( DownstreamStackBusLane[45][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane6_strm0_data          ( DownstreamStackBusLane[45][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane6_strm0_data_valid    ( DownstreamStackBusLane[45][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane6_strm1_ready         ( DownstreamStackBusLane[45][6].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane6_strm1_cntl          ( DownstreamStackBusLane[45][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane6_strm1_data          ( DownstreamStackBusLane[45][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane6_strm1_data_valid    ( DownstreamStackBusLane[45][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane7_strm0_ready         ( DownstreamStackBusLane[45][7].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane7_strm0_cntl          ( DownstreamStackBusLane[45][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane7_strm0_data          ( DownstreamStackBusLane[45][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane7_strm0_data_valid    ( DownstreamStackBusLane[45][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane7_strm1_ready         ( DownstreamStackBusLane[45][7].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane7_strm1_cntl          ( DownstreamStackBusLane[45][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane7_strm1_data          ( DownstreamStackBusLane[45][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane7_strm1_data_valid    ( DownstreamStackBusLane[45][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane8_strm0_ready         ( DownstreamStackBusLane[45][8].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane8_strm0_cntl          ( DownstreamStackBusLane[45][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane8_strm0_data          ( DownstreamStackBusLane[45][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane8_strm0_data_valid    ( DownstreamStackBusLane[45][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane8_strm1_ready         ( DownstreamStackBusLane[45][8].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane8_strm1_cntl          ( DownstreamStackBusLane[45][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane8_strm1_data          ( DownstreamStackBusLane[45][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane8_strm1_data_valid    ( DownstreamStackBusLane[45][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane9_strm0_ready         ( DownstreamStackBusLane[45][9].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane9_strm0_cntl          ( DownstreamStackBusLane[45][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane9_strm0_data          ( DownstreamStackBusLane[45][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane9_strm0_data_valid    ( DownstreamStackBusLane[45][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane9_strm1_ready         ( DownstreamStackBusLane[45][9].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane9_strm1_cntl          ( DownstreamStackBusLane[45][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane9_strm1_data          ( DownstreamStackBusLane[45][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane9_strm1_data_valid    ( DownstreamStackBusLane[45][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane10_strm0_ready         ( DownstreamStackBusLane[45][10].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane10_strm0_cntl          ( DownstreamStackBusLane[45][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane10_strm0_data          ( DownstreamStackBusLane[45][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane10_strm0_data_valid    ( DownstreamStackBusLane[45][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane10_strm1_ready         ( DownstreamStackBusLane[45][10].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane10_strm1_cntl          ( DownstreamStackBusLane[45][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane10_strm1_data          ( DownstreamStackBusLane[45][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane10_strm1_data_valid    ( DownstreamStackBusLane[45][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane11_strm0_ready         ( DownstreamStackBusLane[45][11].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane11_strm0_cntl          ( DownstreamStackBusLane[45][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane11_strm0_data          ( DownstreamStackBusLane[45][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane11_strm0_data_valid    ( DownstreamStackBusLane[45][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane11_strm1_ready         ( DownstreamStackBusLane[45][11].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane11_strm1_cntl          ( DownstreamStackBusLane[45][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane11_strm1_data          ( DownstreamStackBusLane[45][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane11_strm1_data_valid    ( DownstreamStackBusLane[45][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane12_strm0_ready         ( DownstreamStackBusLane[45][12].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane12_strm0_cntl          ( DownstreamStackBusLane[45][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane12_strm0_data          ( DownstreamStackBusLane[45][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane12_strm0_data_valid    ( DownstreamStackBusLane[45][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane12_strm1_ready         ( DownstreamStackBusLane[45][12].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane12_strm1_cntl          ( DownstreamStackBusLane[45][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane12_strm1_data          ( DownstreamStackBusLane[45][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane12_strm1_data_valid    ( DownstreamStackBusLane[45][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane13_strm0_ready         ( DownstreamStackBusLane[45][13].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane13_strm0_cntl          ( DownstreamStackBusLane[45][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane13_strm0_data          ( DownstreamStackBusLane[45][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane13_strm0_data_valid    ( DownstreamStackBusLane[45][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane13_strm1_ready         ( DownstreamStackBusLane[45][13].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane13_strm1_cntl          ( DownstreamStackBusLane[45][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane13_strm1_data          ( DownstreamStackBusLane[45][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane13_strm1_data_valid    ( DownstreamStackBusLane[45][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane14_strm0_ready         ( DownstreamStackBusLane[45][14].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane14_strm0_cntl          ( DownstreamStackBusLane[45][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane14_strm0_data          ( DownstreamStackBusLane[45][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane14_strm0_data_valid    ( DownstreamStackBusLane[45][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane14_strm1_ready         ( DownstreamStackBusLane[45][14].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane14_strm1_cntl          ( DownstreamStackBusLane[45][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane14_strm1_data          ( DownstreamStackBusLane[45][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane14_strm1_data_valid    ( DownstreamStackBusLane[45][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane15_strm0_ready         ( DownstreamStackBusLane[45][15].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane15_strm0_cntl          ( DownstreamStackBusLane[45][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane15_strm0_data          ( DownstreamStackBusLane[45][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane15_strm0_data_valid    ( DownstreamStackBusLane[45][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane15_strm1_ready         ( DownstreamStackBusLane[45][15].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane15_strm1_cntl          ( DownstreamStackBusLane[45][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane15_strm1_data          ( DownstreamStackBusLane[45][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane15_strm1_data_valid    ( DownstreamStackBusLane[45][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane16_strm0_ready         ( DownstreamStackBusLane[45][16].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane16_strm0_cntl          ( DownstreamStackBusLane[45][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane16_strm0_data          ( DownstreamStackBusLane[45][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane16_strm0_data_valid    ( DownstreamStackBusLane[45][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane16_strm1_ready         ( DownstreamStackBusLane[45][16].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane16_strm1_cntl          ( DownstreamStackBusLane[45][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane16_strm1_data          ( DownstreamStackBusLane[45][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane16_strm1_data_valid    ( DownstreamStackBusLane[45][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane17_strm0_ready         ( DownstreamStackBusLane[45][17].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane17_strm0_cntl          ( DownstreamStackBusLane[45][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane17_strm0_data          ( DownstreamStackBusLane[45][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane17_strm0_data_valid    ( DownstreamStackBusLane[45][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane17_strm1_ready         ( DownstreamStackBusLane[45][17].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane17_strm1_cntl          ( DownstreamStackBusLane[45][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane17_strm1_data          ( DownstreamStackBusLane[45][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane17_strm1_data_valid    ( DownstreamStackBusLane[45][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane18_strm0_ready         ( DownstreamStackBusLane[45][18].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane18_strm0_cntl          ( DownstreamStackBusLane[45][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane18_strm0_data          ( DownstreamStackBusLane[45][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane18_strm0_data_valid    ( DownstreamStackBusLane[45][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane18_strm1_ready         ( DownstreamStackBusLane[45][18].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane18_strm1_cntl          ( DownstreamStackBusLane[45][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane18_strm1_data          ( DownstreamStackBusLane[45][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane18_strm1_data_valid    ( DownstreamStackBusLane[45][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane19_strm0_ready         ( DownstreamStackBusLane[45][19].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane19_strm0_cntl          ( DownstreamStackBusLane[45][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane19_strm0_data          ( DownstreamStackBusLane[45][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane19_strm0_data_valid    ( DownstreamStackBusLane[45][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane19_strm1_ready         ( DownstreamStackBusLane[45][19].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane19_strm1_cntl          ( DownstreamStackBusLane[45][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane19_strm1_data          ( DownstreamStackBusLane[45][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane19_strm1_data_valid    ( DownstreamStackBusLane[45][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane20_strm0_ready         ( DownstreamStackBusLane[45][20].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane20_strm0_cntl          ( DownstreamStackBusLane[45][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane20_strm0_data          ( DownstreamStackBusLane[45][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane20_strm0_data_valid    ( DownstreamStackBusLane[45][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane20_strm1_ready         ( DownstreamStackBusLane[45][20].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane20_strm1_cntl          ( DownstreamStackBusLane[45][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane20_strm1_data          ( DownstreamStackBusLane[45][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane20_strm1_data_valid    ( DownstreamStackBusLane[45][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane21_strm0_ready         ( DownstreamStackBusLane[45][21].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane21_strm0_cntl          ( DownstreamStackBusLane[45][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane21_strm0_data          ( DownstreamStackBusLane[45][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane21_strm0_data_valid    ( DownstreamStackBusLane[45][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane21_strm1_ready         ( DownstreamStackBusLane[45][21].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane21_strm1_cntl          ( DownstreamStackBusLane[45][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane21_strm1_data          ( DownstreamStackBusLane[45][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane21_strm1_data_valid    ( DownstreamStackBusLane[45][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane22_strm0_ready         ( DownstreamStackBusLane[45][22].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane22_strm0_cntl          ( DownstreamStackBusLane[45][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane22_strm0_data          ( DownstreamStackBusLane[45][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane22_strm0_data_valid    ( DownstreamStackBusLane[45][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane22_strm1_ready         ( DownstreamStackBusLane[45][22].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane22_strm1_cntl          ( DownstreamStackBusLane[45][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane22_strm1_data          ( DownstreamStackBusLane[45][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane22_strm1_data_valid    ( DownstreamStackBusLane[45][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane23_strm0_ready         ( DownstreamStackBusLane[45][23].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane23_strm0_cntl          ( DownstreamStackBusLane[45][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane23_strm0_data          ( DownstreamStackBusLane[45][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane23_strm0_data_valid    ( DownstreamStackBusLane[45][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane23_strm1_ready         ( DownstreamStackBusLane[45][23].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane23_strm1_cntl          ( DownstreamStackBusLane[45][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane23_strm1_data          ( DownstreamStackBusLane[45][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane23_strm1_data_valid    ( DownstreamStackBusLane[45][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane24_strm0_ready         ( DownstreamStackBusLane[45][24].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane24_strm0_cntl          ( DownstreamStackBusLane[45][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane24_strm0_data          ( DownstreamStackBusLane[45][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane24_strm0_data_valid    ( DownstreamStackBusLane[45][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane24_strm1_ready         ( DownstreamStackBusLane[45][24].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane24_strm1_cntl          ( DownstreamStackBusLane[45][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane24_strm1_data          ( DownstreamStackBusLane[45][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane24_strm1_data_valid    ( DownstreamStackBusLane[45][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane25_strm0_ready         ( DownstreamStackBusLane[45][25].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane25_strm0_cntl          ( DownstreamStackBusLane[45][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane25_strm0_data          ( DownstreamStackBusLane[45][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane25_strm0_data_valid    ( DownstreamStackBusLane[45][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane25_strm1_ready         ( DownstreamStackBusLane[45][25].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane25_strm1_cntl          ( DownstreamStackBusLane[45][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane25_strm1_data          ( DownstreamStackBusLane[45][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane25_strm1_data_valid    ( DownstreamStackBusLane[45][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane26_strm0_ready         ( DownstreamStackBusLane[45][26].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane26_strm0_cntl          ( DownstreamStackBusLane[45][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane26_strm0_data          ( DownstreamStackBusLane[45][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane26_strm0_data_valid    ( DownstreamStackBusLane[45][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane26_strm1_ready         ( DownstreamStackBusLane[45][26].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane26_strm1_cntl          ( DownstreamStackBusLane[45][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane26_strm1_data          ( DownstreamStackBusLane[45][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane26_strm1_data_valid    ( DownstreamStackBusLane[45][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane27_strm0_ready         ( DownstreamStackBusLane[45][27].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane27_strm0_cntl          ( DownstreamStackBusLane[45][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane27_strm0_data          ( DownstreamStackBusLane[45][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane27_strm0_data_valid    ( DownstreamStackBusLane[45][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane27_strm1_ready         ( DownstreamStackBusLane[45][27].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane27_strm1_cntl          ( DownstreamStackBusLane[45][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane27_strm1_data          ( DownstreamStackBusLane[45][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane27_strm1_data_valid    ( DownstreamStackBusLane[45][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane28_strm0_ready         ( DownstreamStackBusLane[45][28].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane28_strm0_cntl          ( DownstreamStackBusLane[45][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane28_strm0_data          ( DownstreamStackBusLane[45][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane28_strm0_data_valid    ( DownstreamStackBusLane[45][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane28_strm1_ready         ( DownstreamStackBusLane[45][28].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane28_strm1_cntl          ( DownstreamStackBusLane[45][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane28_strm1_data          ( DownstreamStackBusLane[45][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane28_strm1_data_valid    ( DownstreamStackBusLane[45][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane29_strm0_ready         ( DownstreamStackBusLane[45][29].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane29_strm0_cntl          ( DownstreamStackBusLane[45][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane29_strm0_data          ( DownstreamStackBusLane[45][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane29_strm0_data_valid    ( DownstreamStackBusLane[45][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane29_strm1_ready         ( DownstreamStackBusLane[45][29].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane29_strm1_cntl          ( DownstreamStackBusLane[45][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane29_strm1_data          ( DownstreamStackBusLane[45][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane29_strm1_data_valid    ( DownstreamStackBusLane[45][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane30_strm0_ready         ( DownstreamStackBusLane[45][30].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane30_strm0_cntl          ( DownstreamStackBusLane[45][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane30_strm0_data          ( DownstreamStackBusLane[45][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane30_strm0_data_valid    ( DownstreamStackBusLane[45][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane30_strm1_ready         ( DownstreamStackBusLane[45][30].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane30_strm1_cntl          ( DownstreamStackBusLane[45][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane30_strm1_data          ( DownstreamStackBusLane[45][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane30_strm1_data_valid    ( DownstreamStackBusLane[45][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 45, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane31_strm0_ready         ( DownstreamStackBusLane[45][31].pe__std__lane_strm0_ready              ),      
        .std__pe45__lane31_strm0_cntl          ( DownstreamStackBusLane[45][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe45__lane31_strm0_data          ( DownstreamStackBusLane[45][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe45__lane31_strm0_data_valid    ( DownstreamStackBusLane[45][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__std__lane31_strm1_ready         ( DownstreamStackBusLane[45][31].pe__std__lane_strm1_ready              ),      
        .std__pe45__lane31_strm1_cntl          ( DownstreamStackBusLane[45][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe45__lane31_strm1_data          ( DownstreamStackBusLane[45][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe45__lane31_strm1_data_valid    ( DownstreamStackBusLane[45][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane0_strm0_ready         ( DownstreamStackBusLane[46][0].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane0_strm0_cntl          ( DownstreamStackBusLane[46][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane0_strm0_data          ( DownstreamStackBusLane[46][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane0_strm0_data_valid    ( DownstreamStackBusLane[46][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane0_strm1_ready         ( DownstreamStackBusLane[46][0].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane0_strm1_cntl          ( DownstreamStackBusLane[46][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane0_strm1_data          ( DownstreamStackBusLane[46][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane0_strm1_data_valid    ( DownstreamStackBusLane[46][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane1_strm0_ready         ( DownstreamStackBusLane[46][1].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane1_strm0_cntl          ( DownstreamStackBusLane[46][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane1_strm0_data          ( DownstreamStackBusLane[46][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane1_strm0_data_valid    ( DownstreamStackBusLane[46][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane1_strm1_ready         ( DownstreamStackBusLane[46][1].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane1_strm1_cntl          ( DownstreamStackBusLane[46][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane1_strm1_data          ( DownstreamStackBusLane[46][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane1_strm1_data_valid    ( DownstreamStackBusLane[46][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane2_strm0_ready         ( DownstreamStackBusLane[46][2].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane2_strm0_cntl          ( DownstreamStackBusLane[46][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane2_strm0_data          ( DownstreamStackBusLane[46][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane2_strm0_data_valid    ( DownstreamStackBusLane[46][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane2_strm1_ready         ( DownstreamStackBusLane[46][2].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane2_strm1_cntl          ( DownstreamStackBusLane[46][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane2_strm1_data          ( DownstreamStackBusLane[46][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane2_strm1_data_valid    ( DownstreamStackBusLane[46][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane3_strm0_ready         ( DownstreamStackBusLane[46][3].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane3_strm0_cntl          ( DownstreamStackBusLane[46][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane3_strm0_data          ( DownstreamStackBusLane[46][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane3_strm0_data_valid    ( DownstreamStackBusLane[46][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane3_strm1_ready         ( DownstreamStackBusLane[46][3].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane3_strm1_cntl          ( DownstreamStackBusLane[46][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane3_strm1_data          ( DownstreamStackBusLane[46][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane3_strm1_data_valid    ( DownstreamStackBusLane[46][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane4_strm0_ready         ( DownstreamStackBusLane[46][4].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane4_strm0_cntl          ( DownstreamStackBusLane[46][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane4_strm0_data          ( DownstreamStackBusLane[46][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane4_strm0_data_valid    ( DownstreamStackBusLane[46][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane4_strm1_ready         ( DownstreamStackBusLane[46][4].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane4_strm1_cntl          ( DownstreamStackBusLane[46][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane4_strm1_data          ( DownstreamStackBusLane[46][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane4_strm1_data_valid    ( DownstreamStackBusLane[46][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane5_strm0_ready         ( DownstreamStackBusLane[46][5].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane5_strm0_cntl          ( DownstreamStackBusLane[46][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane5_strm0_data          ( DownstreamStackBusLane[46][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane5_strm0_data_valid    ( DownstreamStackBusLane[46][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane5_strm1_ready         ( DownstreamStackBusLane[46][5].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane5_strm1_cntl          ( DownstreamStackBusLane[46][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane5_strm1_data          ( DownstreamStackBusLane[46][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane5_strm1_data_valid    ( DownstreamStackBusLane[46][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane6_strm0_ready         ( DownstreamStackBusLane[46][6].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane6_strm0_cntl          ( DownstreamStackBusLane[46][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane6_strm0_data          ( DownstreamStackBusLane[46][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane6_strm0_data_valid    ( DownstreamStackBusLane[46][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane6_strm1_ready         ( DownstreamStackBusLane[46][6].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane6_strm1_cntl          ( DownstreamStackBusLane[46][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane6_strm1_data          ( DownstreamStackBusLane[46][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane6_strm1_data_valid    ( DownstreamStackBusLane[46][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane7_strm0_ready         ( DownstreamStackBusLane[46][7].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane7_strm0_cntl          ( DownstreamStackBusLane[46][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane7_strm0_data          ( DownstreamStackBusLane[46][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane7_strm0_data_valid    ( DownstreamStackBusLane[46][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane7_strm1_ready         ( DownstreamStackBusLane[46][7].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane7_strm1_cntl          ( DownstreamStackBusLane[46][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane7_strm1_data          ( DownstreamStackBusLane[46][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane7_strm1_data_valid    ( DownstreamStackBusLane[46][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane8_strm0_ready         ( DownstreamStackBusLane[46][8].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane8_strm0_cntl          ( DownstreamStackBusLane[46][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane8_strm0_data          ( DownstreamStackBusLane[46][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane8_strm0_data_valid    ( DownstreamStackBusLane[46][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane8_strm1_ready         ( DownstreamStackBusLane[46][8].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane8_strm1_cntl          ( DownstreamStackBusLane[46][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane8_strm1_data          ( DownstreamStackBusLane[46][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane8_strm1_data_valid    ( DownstreamStackBusLane[46][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane9_strm0_ready         ( DownstreamStackBusLane[46][9].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane9_strm0_cntl          ( DownstreamStackBusLane[46][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane9_strm0_data          ( DownstreamStackBusLane[46][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane9_strm0_data_valid    ( DownstreamStackBusLane[46][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane9_strm1_ready         ( DownstreamStackBusLane[46][9].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane9_strm1_cntl          ( DownstreamStackBusLane[46][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane9_strm1_data          ( DownstreamStackBusLane[46][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane9_strm1_data_valid    ( DownstreamStackBusLane[46][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane10_strm0_ready         ( DownstreamStackBusLane[46][10].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane10_strm0_cntl          ( DownstreamStackBusLane[46][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane10_strm0_data          ( DownstreamStackBusLane[46][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane10_strm0_data_valid    ( DownstreamStackBusLane[46][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane10_strm1_ready         ( DownstreamStackBusLane[46][10].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane10_strm1_cntl          ( DownstreamStackBusLane[46][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane10_strm1_data          ( DownstreamStackBusLane[46][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane10_strm1_data_valid    ( DownstreamStackBusLane[46][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane11_strm0_ready         ( DownstreamStackBusLane[46][11].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane11_strm0_cntl          ( DownstreamStackBusLane[46][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane11_strm0_data          ( DownstreamStackBusLane[46][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane11_strm0_data_valid    ( DownstreamStackBusLane[46][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane11_strm1_ready         ( DownstreamStackBusLane[46][11].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane11_strm1_cntl          ( DownstreamStackBusLane[46][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane11_strm1_data          ( DownstreamStackBusLane[46][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane11_strm1_data_valid    ( DownstreamStackBusLane[46][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane12_strm0_ready         ( DownstreamStackBusLane[46][12].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane12_strm0_cntl          ( DownstreamStackBusLane[46][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane12_strm0_data          ( DownstreamStackBusLane[46][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane12_strm0_data_valid    ( DownstreamStackBusLane[46][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane12_strm1_ready         ( DownstreamStackBusLane[46][12].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane12_strm1_cntl          ( DownstreamStackBusLane[46][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane12_strm1_data          ( DownstreamStackBusLane[46][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane12_strm1_data_valid    ( DownstreamStackBusLane[46][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane13_strm0_ready         ( DownstreamStackBusLane[46][13].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane13_strm0_cntl          ( DownstreamStackBusLane[46][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane13_strm0_data          ( DownstreamStackBusLane[46][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane13_strm0_data_valid    ( DownstreamStackBusLane[46][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane13_strm1_ready         ( DownstreamStackBusLane[46][13].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane13_strm1_cntl          ( DownstreamStackBusLane[46][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane13_strm1_data          ( DownstreamStackBusLane[46][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane13_strm1_data_valid    ( DownstreamStackBusLane[46][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane14_strm0_ready         ( DownstreamStackBusLane[46][14].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane14_strm0_cntl          ( DownstreamStackBusLane[46][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane14_strm0_data          ( DownstreamStackBusLane[46][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane14_strm0_data_valid    ( DownstreamStackBusLane[46][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane14_strm1_ready         ( DownstreamStackBusLane[46][14].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane14_strm1_cntl          ( DownstreamStackBusLane[46][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane14_strm1_data          ( DownstreamStackBusLane[46][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane14_strm1_data_valid    ( DownstreamStackBusLane[46][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane15_strm0_ready         ( DownstreamStackBusLane[46][15].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane15_strm0_cntl          ( DownstreamStackBusLane[46][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane15_strm0_data          ( DownstreamStackBusLane[46][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane15_strm0_data_valid    ( DownstreamStackBusLane[46][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane15_strm1_ready         ( DownstreamStackBusLane[46][15].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane15_strm1_cntl          ( DownstreamStackBusLane[46][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane15_strm1_data          ( DownstreamStackBusLane[46][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane15_strm1_data_valid    ( DownstreamStackBusLane[46][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane16_strm0_ready         ( DownstreamStackBusLane[46][16].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane16_strm0_cntl          ( DownstreamStackBusLane[46][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane16_strm0_data          ( DownstreamStackBusLane[46][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane16_strm0_data_valid    ( DownstreamStackBusLane[46][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane16_strm1_ready         ( DownstreamStackBusLane[46][16].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane16_strm1_cntl          ( DownstreamStackBusLane[46][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane16_strm1_data          ( DownstreamStackBusLane[46][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane16_strm1_data_valid    ( DownstreamStackBusLane[46][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane17_strm0_ready         ( DownstreamStackBusLane[46][17].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane17_strm0_cntl          ( DownstreamStackBusLane[46][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane17_strm0_data          ( DownstreamStackBusLane[46][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane17_strm0_data_valid    ( DownstreamStackBusLane[46][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane17_strm1_ready         ( DownstreamStackBusLane[46][17].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane17_strm1_cntl          ( DownstreamStackBusLane[46][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane17_strm1_data          ( DownstreamStackBusLane[46][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane17_strm1_data_valid    ( DownstreamStackBusLane[46][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane18_strm0_ready         ( DownstreamStackBusLane[46][18].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane18_strm0_cntl          ( DownstreamStackBusLane[46][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane18_strm0_data          ( DownstreamStackBusLane[46][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane18_strm0_data_valid    ( DownstreamStackBusLane[46][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane18_strm1_ready         ( DownstreamStackBusLane[46][18].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane18_strm1_cntl          ( DownstreamStackBusLane[46][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane18_strm1_data          ( DownstreamStackBusLane[46][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane18_strm1_data_valid    ( DownstreamStackBusLane[46][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane19_strm0_ready         ( DownstreamStackBusLane[46][19].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane19_strm0_cntl          ( DownstreamStackBusLane[46][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane19_strm0_data          ( DownstreamStackBusLane[46][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane19_strm0_data_valid    ( DownstreamStackBusLane[46][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane19_strm1_ready         ( DownstreamStackBusLane[46][19].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane19_strm1_cntl          ( DownstreamStackBusLane[46][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane19_strm1_data          ( DownstreamStackBusLane[46][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane19_strm1_data_valid    ( DownstreamStackBusLane[46][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane20_strm0_ready         ( DownstreamStackBusLane[46][20].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane20_strm0_cntl          ( DownstreamStackBusLane[46][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane20_strm0_data          ( DownstreamStackBusLane[46][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane20_strm0_data_valid    ( DownstreamStackBusLane[46][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane20_strm1_ready         ( DownstreamStackBusLane[46][20].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane20_strm1_cntl          ( DownstreamStackBusLane[46][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane20_strm1_data          ( DownstreamStackBusLane[46][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane20_strm1_data_valid    ( DownstreamStackBusLane[46][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane21_strm0_ready         ( DownstreamStackBusLane[46][21].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane21_strm0_cntl          ( DownstreamStackBusLane[46][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane21_strm0_data          ( DownstreamStackBusLane[46][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane21_strm0_data_valid    ( DownstreamStackBusLane[46][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane21_strm1_ready         ( DownstreamStackBusLane[46][21].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane21_strm1_cntl          ( DownstreamStackBusLane[46][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane21_strm1_data          ( DownstreamStackBusLane[46][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane21_strm1_data_valid    ( DownstreamStackBusLane[46][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane22_strm0_ready         ( DownstreamStackBusLane[46][22].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane22_strm0_cntl          ( DownstreamStackBusLane[46][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane22_strm0_data          ( DownstreamStackBusLane[46][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane22_strm0_data_valid    ( DownstreamStackBusLane[46][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane22_strm1_ready         ( DownstreamStackBusLane[46][22].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane22_strm1_cntl          ( DownstreamStackBusLane[46][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane22_strm1_data          ( DownstreamStackBusLane[46][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane22_strm1_data_valid    ( DownstreamStackBusLane[46][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane23_strm0_ready         ( DownstreamStackBusLane[46][23].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane23_strm0_cntl          ( DownstreamStackBusLane[46][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane23_strm0_data          ( DownstreamStackBusLane[46][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane23_strm0_data_valid    ( DownstreamStackBusLane[46][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane23_strm1_ready         ( DownstreamStackBusLane[46][23].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane23_strm1_cntl          ( DownstreamStackBusLane[46][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane23_strm1_data          ( DownstreamStackBusLane[46][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane23_strm1_data_valid    ( DownstreamStackBusLane[46][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane24_strm0_ready         ( DownstreamStackBusLane[46][24].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane24_strm0_cntl          ( DownstreamStackBusLane[46][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane24_strm0_data          ( DownstreamStackBusLane[46][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane24_strm0_data_valid    ( DownstreamStackBusLane[46][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane24_strm1_ready         ( DownstreamStackBusLane[46][24].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane24_strm1_cntl          ( DownstreamStackBusLane[46][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane24_strm1_data          ( DownstreamStackBusLane[46][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane24_strm1_data_valid    ( DownstreamStackBusLane[46][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane25_strm0_ready         ( DownstreamStackBusLane[46][25].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane25_strm0_cntl          ( DownstreamStackBusLane[46][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane25_strm0_data          ( DownstreamStackBusLane[46][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane25_strm0_data_valid    ( DownstreamStackBusLane[46][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane25_strm1_ready         ( DownstreamStackBusLane[46][25].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane25_strm1_cntl          ( DownstreamStackBusLane[46][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane25_strm1_data          ( DownstreamStackBusLane[46][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane25_strm1_data_valid    ( DownstreamStackBusLane[46][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane26_strm0_ready         ( DownstreamStackBusLane[46][26].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane26_strm0_cntl          ( DownstreamStackBusLane[46][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane26_strm0_data          ( DownstreamStackBusLane[46][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane26_strm0_data_valid    ( DownstreamStackBusLane[46][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane26_strm1_ready         ( DownstreamStackBusLane[46][26].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane26_strm1_cntl          ( DownstreamStackBusLane[46][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane26_strm1_data          ( DownstreamStackBusLane[46][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane26_strm1_data_valid    ( DownstreamStackBusLane[46][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane27_strm0_ready         ( DownstreamStackBusLane[46][27].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane27_strm0_cntl          ( DownstreamStackBusLane[46][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane27_strm0_data          ( DownstreamStackBusLane[46][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane27_strm0_data_valid    ( DownstreamStackBusLane[46][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane27_strm1_ready         ( DownstreamStackBusLane[46][27].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane27_strm1_cntl          ( DownstreamStackBusLane[46][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane27_strm1_data          ( DownstreamStackBusLane[46][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane27_strm1_data_valid    ( DownstreamStackBusLane[46][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane28_strm0_ready         ( DownstreamStackBusLane[46][28].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane28_strm0_cntl          ( DownstreamStackBusLane[46][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane28_strm0_data          ( DownstreamStackBusLane[46][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane28_strm0_data_valid    ( DownstreamStackBusLane[46][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane28_strm1_ready         ( DownstreamStackBusLane[46][28].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane28_strm1_cntl          ( DownstreamStackBusLane[46][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane28_strm1_data          ( DownstreamStackBusLane[46][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane28_strm1_data_valid    ( DownstreamStackBusLane[46][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane29_strm0_ready         ( DownstreamStackBusLane[46][29].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane29_strm0_cntl          ( DownstreamStackBusLane[46][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane29_strm0_data          ( DownstreamStackBusLane[46][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane29_strm0_data_valid    ( DownstreamStackBusLane[46][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane29_strm1_ready         ( DownstreamStackBusLane[46][29].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane29_strm1_cntl          ( DownstreamStackBusLane[46][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane29_strm1_data          ( DownstreamStackBusLane[46][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane29_strm1_data_valid    ( DownstreamStackBusLane[46][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane30_strm0_ready         ( DownstreamStackBusLane[46][30].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane30_strm0_cntl          ( DownstreamStackBusLane[46][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane30_strm0_data          ( DownstreamStackBusLane[46][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane30_strm0_data_valid    ( DownstreamStackBusLane[46][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane30_strm1_ready         ( DownstreamStackBusLane[46][30].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane30_strm1_cntl          ( DownstreamStackBusLane[46][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane30_strm1_data          ( DownstreamStackBusLane[46][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane30_strm1_data_valid    ( DownstreamStackBusLane[46][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 46, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane31_strm0_ready         ( DownstreamStackBusLane[46][31].pe__std__lane_strm0_ready              ),      
        .std__pe46__lane31_strm0_cntl          ( DownstreamStackBusLane[46][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe46__lane31_strm0_data          ( DownstreamStackBusLane[46][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe46__lane31_strm0_data_valid    ( DownstreamStackBusLane[46][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__std__lane31_strm1_ready         ( DownstreamStackBusLane[46][31].pe__std__lane_strm1_ready              ),      
        .std__pe46__lane31_strm1_cntl          ( DownstreamStackBusLane[46][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe46__lane31_strm1_data          ( DownstreamStackBusLane[46][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe46__lane31_strm1_data_valid    ( DownstreamStackBusLane[46][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane0_strm0_ready         ( DownstreamStackBusLane[47][0].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane0_strm0_cntl          ( DownstreamStackBusLane[47][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane0_strm0_data          ( DownstreamStackBusLane[47][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane0_strm0_data_valid    ( DownstreamStackBusLane[47][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane0_strm1_ready         ( DownstreamStackBusLane[47][0].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane0_strm1_cntl          ( DownstreamStackBusLane[47][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane0_strm1_data          ( DownstreamStackBusLane[47][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane0_strm1_data_valid    ( DownstreamStackBusLane[47][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane1_strm0_ready         ( DownstreamStackBusLane[47][1].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane1_strm0_cntl          ( DownstreamStackBusLane[47][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane1_strm0_data          ( DownstreamStackBusLane[47][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane1_strm0_data_valid    ( DownstreamStackBusLane[47][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane1_strm1_ready         ( DownstreamStackBusLane[47][1].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane1_strm1_cntl          ( DownstreamStackBusLane[47][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane1_strm1_data          ( DownstreamStackBusLane[47][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane1_strm1_data_valid    ( DownstreamStackBusLane[47][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane2_strm0_ready         ( DownstreamStackBusLane[47][2].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane2_strm0_cntl          ( DownstreamStackBusLane[47][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane2_strm0_data          ( DownstreamStackBusLane[47][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane2_strm0_data_valid    ( DownstreamStackBusLane[47][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane2_strm1_ready         ( DownstreamStackBusLane[47][2].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane2_strm1_cntl          ( DownstreamStackBusLane[47][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane2_strm1_data          ( DownstreamStackBusLane[47][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane2_strm1_data_valid    ( DownstreamStackBusLane[47][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane3_strm0_ready         ( DownstreamStackBusLane[47][3].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane3_strm0_cntl          ( DownstreamStackBusLane[47][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane3_strm0_data          ( DownstreamStackBusLane[47][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane3_strm0_data_valid    ( DownstreamStackBusLane[47][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane3_strm1_ready         ( DownstreamStackBusLane[47][3].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane3_strm1_cntl          ( DownstreamStackBusLane[47][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane3_strm1_data          ( DownstreamStackBusLane[47][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane3_strm1_data_valid    ( DownstreamStackBusLane[47][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane4_strm0_ready         ( DownstreamStackBusLane[47][4].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane4_strm0_cntl          ( DownstreamStackBusLane[47][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane4_strm0_data          ( DownstreamStackBusLane[47][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane4_strm0_data_valid    ( DownstreamStackBusLane[47][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane4_strm1_ready         ( DownstreamStackBusLane[47][4].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane4_strm1_cntl          ( DownstreamStackBusLane[47][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane4_strm1_data          ( DownstreamStackBusLane[47][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane4_strm1_data_valid    ( DownstreamStackBusLane[47][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane5_strm0_ready         ( DownstreamStackBusLane[47][5].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane5_strm0_cntl          ( DownstreamStackBusLane[47][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane5_strm0_data          ( DownstreamStackBusLane[47][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane5_strm0_data_valid    ( DownstreamStackBusLane[47][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane5_strm1_ready         ( DownstreamStackBusLane[47][5].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane5_strm1_cntl          ( DownstreamStackBusLane[47][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane5_strm1_data          ( DownstreamStackBusLane[47][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane5_strm1_data_valid    ( DownstreamStackBusLane[47][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane6_strm0_ready         ( DownstreamStackBusLane[47][6].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane6_strm0_cntl          ( DownstreamStackBusLane[47][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane6_strm0_data          ( DownstreamStackBusLane[47][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane6_strm0_data_valid    ( DownstreamStackBusLane[47][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane6_strm1_ready         ( DownstreamStackBusLane[47][6].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane6_strm1_cntl          ( DownstreamStackBusLane[47][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane6_strm1_data          ( DownstreamStackBusLane[47][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane6_strm1_data_valid    ( DownstreamStackBusLane[47][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane7_strm0_ready         ( DownstreamStackBusLane[47][7].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane7_strm0_cntl          ( DownstreamStackBusLane[47][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane7_strm0_data          ( DownstreamStackBusLane[47][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane7_strm0_data_valid    ( DownstreamStackBusLane[47][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane7_strm1_ready         ( DownstreamStackBusLane[47][7].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane7_strm1_cntl          ( DownstreamStackBusLane[47][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane7_strm1_data          ( DownstreamStackBusLane[47][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane7_strm1_data_valid    ( DownstreamStackBusLane[47][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane8_strm0_ready         ( DownstreamStackBusLane[47][8].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane8_strm0_cntl          ( DownstreamStackBusLane[47][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane8_strm0_data          ( DownstreamStackBusLane[47][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane8_strm0_data_valid    ( DownstreamStackBusLane[47][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane8_strm1_ready         ( DownstreamStackBusLane[47][8].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane8_strm1_cntl          ( DownstreamStackBusLane[47][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane8_strm1_data          ( DownstreamStackBusLane[47][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane8_strm1_data_valid    ( DownstreamStackBusLane[47][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane9_strm0_ready         ( DownstreamStackBusLane[47][9].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane9_strm0_cntl          ( DownstreamStackBusLane[47][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane9_strm0_data          ( DownstreamStackBusLane[47][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane9_strm0_data_valid    ( DownstreamStackBusLane[47][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane9_strm1_ready         ( DownstreamStackBusLane[47][9].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane9_strm1_cntl          ( DownstreamStackBusLane[47][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane9_strm1_data          ( DownstreamStackBusLane[47][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane9_strm1_data_valid    ( DownstreamStackBusLane[47][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane10_strm0_ready         ( DownstreamStackBusLane[47][10].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane10_strm0_cntl          ( DownstreamStackBusLane[47][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane10_strm0_data          ( DownstreamStackBusLane[47][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane10_strm0_data_valid    ( DownstreamStackBusLane[47][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane10_strm1_ready         ( DownstreamStackBusLane[47][10].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane10_strm1_cntl          ( DownstreamStackBusLane[47][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane10_strm1_data          ( DownstreamStackBusLane[47][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane10_strm1_data_valid    ( DownstreamStackBusLane[47][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane11_strm0_ready         ( DownstreamStackBusLane[47][11].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane11_strm0_cntl          ( DownstreamStackBusLane[47][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane11_strm0_data          ( DownstreamStackBusLane[47][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane11_strm0_data_valid    ( DownstreamStackBusLane[47][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane11_strm1_ready         ( DownstreamStackBusLane[47][11].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane11_strm1_cntl          ( DownstreamStackBusLane[47][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane11_strm1_data          ( DownstreamStackBusLane[47][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane11_strm1_data_valid    ( DownstreamStackBusLane[47][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane12_strm0_ready         ( DownstreamStackBusLane[47][12].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane12_strm0_cntl          ( DownstreamStackBusLane[47][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane12_strm0_data          ( DownstreamStackBusLane[47][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane12_strm0_data_valid    ( DownstreamStackBusLane[47][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane12_strm1_ready         ( DownstreamStackBusLane[47][12].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane12_strm1_cntl          ( DownstreamStackBusLane[47][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane12_strm1_data          ( DownstreamStackBusLane[47][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane12_strm1_data_valid    ( DownstreamStackBusLane[47][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane13_strm0_ready         ( DownstreamStackBusLane[47][13].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane13_strm0_cntl          ( DownstreamStackBusLane[47][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane13_strm0_data          ( DownstreamStackBusLane[47][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane13_strm0_data_valid    ( DownstreamStackBusLane[47][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane13_strm1_ready         ( DownstreamStackBusLane[47][13].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane13_strm1_cntl          ( DownstreamStackBusLane[47][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane13_strm1_data          ( DownstreamStackBusLane[47][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane13_strm1_data_valid    ( DownstreamStackBusLane[47][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane14_strm0_ready         ( DownstreamStackBusLane[47][14].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane14_strm0_cntl          ( DownstreamStackBusLane[47][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane14_strm0_data          ( DownstreamStackBusLane[47][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane14_strm0_data_valid    ( DownstreamStackBusLane[47][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane14_strm1_ready         ( DownstreamStackBusLane[47][14].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane14_strm1_cntl          ( DownstreamStackBusLane[47][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane14_strm1_data          ( DownstreamStackBusLane[47][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane14_strm1_data_valid    ( DownstreamStackBusLane[47][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane15_strm0_ready         ( DownstreamStackBusLane[47][15].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane15_strm0_cntl          ( DownstreamStackBusLane[47][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane15_strm0_data          ( DownstreamStackBusLane[47][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane15_strm0_data_valid    ( DownstreamStackBusLane[47][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane15_strm1_ready         ( DownstreamStackBusLane[47][15].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane15_strm1_cntl          ( DownstreamStackBusLane[47][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane15_strm1_data          ( DownstreamStackBusLane[47][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane15_strm1_data_valid    ( DownstreamStackBusLane[47][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane16_strm0_ready         ( DownstreamStackBusLane[47][16].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane16_strm0_cntl          ( DownstreamStackBusLane[47][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane16_strm0_data          ( DownstreamStackBusLane[47][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane16_strm0_data_valid    ( DownstreamStackBusLane[47][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane16_strm1_ready         ( DownstreamStackBusLane[47][16].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane16_strm1_cntl          ( DownstreamStackBusLane[47][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane16_strm1_data          ( DownstreamStackBusLane[47][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane16_strm1_data_valid    ( DownstreamStackBusLane[47][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane17_strm0_ready         ( DownstreamStackBusLane[47][17].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane17_strm0_cntl          ( DownstreamStackBusLane[47][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane17_strm0_data          ( DownstreamStackBusLane[47][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane17_strm0_data_valid    ( DownstreamStackBusLane[47][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane17_strm1_ready         ( DownstreamStackBusLane[47][17].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane17_strm1_cntl          ( DownstreamStackBusLane[47][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane17_strm1_data          ( DownstreamStackBusLane[47][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane17_strm1_data_valid    ( DownstreamStackBusLane[47][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane18_strm0_ready         ( DownstreamStackBusLane[47][18].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane18_strm0_cntl          ( DownstreamStackBusLane[47][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane18_strm0_data          ( DownstreamStackBusLane[47][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane18_strm0_data_valid    ( DownstreamStackBusLane[47][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane18_strm1_ready         ( DownstreamStackBusLane[47][18].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane18_strm1_cntl          ( DownstreamStackBusLane[47][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane18_strm1_data          ( DownstreamStackBusLane[47][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane18_strm1_data_valid    ( DownstreamStackBusLane[47][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane19_strm0_ready         ( DownstreamStackBusLane[47][19].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane19_strm0_cntl          ( DownstreamStackBusLane[47][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane19_strm0_data          ( DownstreamStackBusLane[47][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane19_strm0_data_valid    ( DownstreamStackBusLane[47][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane19_strm1_ready         ( DownstreamStackBusLane[47][19].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane19_strm1_cntl          ( DownstreamStackBusLane[47][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane19_strm1_data          ( DownstreamStackBusLane[47][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane19_strm1_data_valid    ( DownstreamStackBusLane[47][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane20_strm0_ready         ( DownstreamStackBusLane[47][20].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane20_strm0_cntl          ( DownstreamStackBusLane[47][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane20_strm0_data          ( DownstreamStackBusLane[47][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane20_strm0_data_valid    ( DownstreamStackBusLane[47][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane20_strm1_ready         ( DownstreamStackBusLane[47][20].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane20_strm1_cntl          ( DownstreamStackBusLane[47][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane20_strm1_data          ( DownstreamStackBusLane[47][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane20_strm1_data_valid    ( DownstreamStackBusLane[47][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane21_strm0_ready         ( DownstreamStackBusLane[47][21].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane21_strm0_cntl          ( DownstreamStackBusLane[47][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane21_strm0_data          ( DownstreamStackBusLane[47][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane21_strm0_data_valid    ( DownstreamStackBusLane[47][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane21_strm1_ready         ( DownstreamStackBusLane[47][21].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane21_strm1_cntl          ( DownstreamStackBusLane[47][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane21_strm1_data          ( DownstreamStackBusLane[47][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane21_strm1_data_valid    ( DownstreamStackBusLane[47][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane22_strm0_ready         ( DownstreamStackBusLane[47][22].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane22_strm0_cntl          ( DownstreamStackBusLane[47][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane22_strm0_data          ( DownstreamStackBusLane[47][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane22_strm0_data_valid    ( DownstreamStackBusLane[47][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane22_strm1_ready         ( DownstreamStackBusLane[47][22].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane22_strm1_cntl          ( DownstreamStackBusLane[47][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane22_strm1_data          ( DownstreamStackBusLane[47][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane22_strm1_data_valid    ( DownstreamStackBusLane[47][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane23_strm0_ready         ( DownstreamStackBusLane[47][23].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane23_strm0_cntl          ( DownstreamStackBusLane[47][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane23_strm0_data          ( DownstreamStackBusLane[47][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane23_strm0_data_valid    ( DownstreamStackBusLane[47][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane23_strm1_ready         ( DownstreamStackBusLane[47][23].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane23_strm1_cntl          ( DownstreamStackBusLane[47][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane23_strm1_data          ( DownstreamStackBusLane[47][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane23_strm1_data_valid    ( DownstreamStackBusLane[47][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane24_strm0_ready         ( DownstreamStackBusLane[47][24].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane24_strm0_cntl          ( DownstreamStackBusLane[47][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane24_strm0_data          ( DownstreamStackBusLane[47][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane24_strm0_data_valid    ( DownstreamStackBusLane[47][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane24_strm1_ready         ( DownstreamStackBusLane[47][24].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane24_strm1_cntl          ( DownstreamStackBusLane[47][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane24_strm1_data          ( DownstreamStackBusLane[47][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane24_strm1_data_valid    ( DownstreamStackBusLane[47][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane25_strm0_ready         ( DownstreamStackBusLane[47][25].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane25_strm0_cntl          ( DownstreamStackBusLane[47][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane25_strm0_data          ( DownstreamStackBusLane[47][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane25_strm0_data_valid    ( DownstreamStackBusLane[47][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane25_strm1_ready         ( DownstreamStackBusLane[47][25].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane25_strm1_cntl          ( DownstreamStackBusLane[47][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane25_strm1_data          ( DownstreamStackBusLane[47][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane25_strm1_data_valid    ( DownstreamStackBusLane[47][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane26_strm0_ready         ( DownstreamStackBusLane[47][26].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane26_strm0_cntl          ( DownstreamStackBusLane[47][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane26_strm0_data          ( DownstreamStackBusLane[47][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane26_strm0_data_valid    ( DownstreamStackBusLane[47][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane26_strm1_ready         ( DownstreamStackBusLane[47][26].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane26_strm1_cntl          ( DownstreamStackBusLane[47][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane26_strm1_data          ( DownstreamStackBusLane[47][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane26_strm1_data_valid    ( DownstreamStackBusLane[47][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane27_strm0_ready         ( DownstreamStackBusLane[47][27].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane27_strm0_cntl          ( DownstreamStackBusLane[47][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane27_strm0_data          ( DownstreamStackBusLane[47][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane27_strm0_data_valid    ( DownstreamStackBusLane[47][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane27_strm1_ready         ( DownstreamStackBusLane[47][27].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane27_strm1_cntl          ( DownstreamStackBusLane[47][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane27_strm1_data          ( DownstreamStackBusLane[47][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane27_strm1_data_valid    ( DownstreamStackBusLane[47][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane28_strm0_ready         ( DownstreamStackBusLane[47][28].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane28_strm0_cntl          ( DownstreamStackBusLane[47][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane28_strm0_data          ( DownstreamStackBusLane[47][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane28_strm0_data_valid    ( DownstreamStackBusLane[47][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane28_strm1_ready         ( DownstreamStackBusLane[47][28].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane28_strm1_cntl          ( DownstreamStackBusLane[47][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane28_strm1_data          ( DownstreamStackBusLane[47][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane28_strm1_data_valid    ( DownstreamStackBusLane[47][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane29_strm0_ready         ( DownstreamStackBusLane[47][29].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane29_strm0_cntl          ( DownstreamStackBusLane[47][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane29_strm0_data          ( DownstreamStackBusLane[47][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane29_strm0_data_valid    ( DownstreamStackBusLane[47][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane29_strm1_ready         ( DownstreamStackBusLane[47][29].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane29_strm1_cntl          ( DownstreamStackBusLane[47][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane29_strm1_data          ( DownstreamStackBusLane[47][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane29_strm1_data_valid    ( DownstreamStackBusLane[47][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane30_strm0_ready         ( DownstreamStackBusLane[47][30].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane30_strm0_cntl          ( DownstreamStackBusLane[47][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane30_strm0_data          ( DownstreamStackBusLane[47][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane30_strm0_data_valid    ( DownstreamStackBusLane[47][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane30_strm1_ready         ( DownstreamStackBusLane[47][30].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane30_strm1_cntl          ( DownstreamStackBusLane[47][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane30_strm1_data          ( DownstreamStackBusLane[47][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane30_strm1_data_valid    ( DownstreamStackBusLane[47][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 47, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane31_strm0_ready         ( DownstreamStackBusLane[47][31].pe__std__lane_strm0_ready              ),      
        .std__pe47__lane31_strm0_cntl          ( DownstreamStackBusLane[47][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe47__lane31_strm0_data          ( DownstreamStackBusLane[47][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe47__lane31_strm0_data_valid    ( DownstreamStackBusLane[47][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__std__lane31_strm1_ready         ( DownstreamStackBusLane[47][31].pe__std__lane_strm1_ready              ),      
        .std__pe47__lane31_strm1_cntl          ( DownstreamStackBusLane[47][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe47__lane31_strm1_data          ( DownstreamStackBusLane[47][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe47__lane31_strm1_data_valid    ( DownstreamStackBusLane[47][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane0_strm0_ready         ( DownstreamStackBusLane[48][0].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane0_strm0_cntl          ( DownstreamStackBusLane[48][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane0_strm0_data          ( DownstreamStackBusLane[48][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane0_strm0_data_valid    ( DownstreamStackBusLane[48][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane0_strm1_ready         ( DownstreamStackBusLane[48][0].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane0_strm1_cntl          ( DownstreamStackBusLane[48][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane0_strm1_data          ( DownstreamStackBusLane[48][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane0_strm1_data_valid    ( DownstreamStackBusLane[48][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane1_strm0_ready         ( DownstreamStackBusLane[48][1].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane1_strm0_cntl          ( DownstreamStackBusLane[48][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane1_strm0_data          ( DownstreamStackBusLane[48][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane1_strm0_data_valid    ( DownstreamStackBusLane[48][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane1_strm1_ready         ( DownstreamStackBusLane[48][1].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane1_strm1_cntl          ( DownstreamStackBusLane[48][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane1_strm1_data          ( DownstreamStackBusLane[48][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane1_strm1_data_valid    ( DownstreamStackBusLane[48][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane2_strm0_ready         ( DownstreamStackBusLane[48][2].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane2_strm0_cntl          ( DownstreamStackBusLane[48][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane2_strm0_data          ( DownstreamStackBusLane[48][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane2_strm0_data_valid    ( DownstreamStackBusLane[48][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane2_strm1_ready         ( DownstreamStackBusLane[48][2].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane2_strm1_cntl          ( DownstreamStackBusLane[48][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane2_strm1_data          ( DownstreamStackBusLane[48][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane2_strm1_data_valid    ( DownstreamStackBusLane[48][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane3_strm0_ready         ( DownstreamStackBusLane[48][3].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane3_strm0_cntl          ( DownstreamStackBusLane[48][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane3_strm0_data          ( DownstreamStackBusLane[48][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane3_strm0_data_valid    ( DownstreamStackBusLane[48][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane3_strm1_ready         ( DownstreamStackBusLane[48][3].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane3_strm1_cntl          ( DownstreamStackBusLane[48][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane3_strm1_data          ( DownstreamStackBusLane[48][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane3_strm1_data_valid    ( DownstreamStackBusLane[48][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane4_strm0_ready         ( DownstreamStackBusLane[48][4].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane4_strm0_cntl          ( DownstreamStackBusLane[48][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane4_strm0_data          ( DownstreamStackBusLane[48][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane4_strm0_data_valid    ( DownstreamStackBusLane[48][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane4_strm1_ready         ( DownstreamStackBusLane[48][4].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane4_strm1_cntl          ( DownstreamStackBusLane[48][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane4_strm1_data          ( DownstreamStackBusLane[48][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane4_strm1_data_valid    ( DownstreamStackBusLane[48][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane5_strm0_ready         ( DownstreamStackBusLane[48][5].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane5_strm0_cntl          ( DownstreamStackBusLane[48][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane5_strm0_data          ( DownstreamStackBusLane[48][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane5_strm0_data_valid    ( DownstreamStackBusLane[48][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane5_strm1_ready         ( DownstreamStackBusLane[48][5].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane5_strm1_cntl          ( DownstreamStackBusLane[48][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane5_strm1_data          ( DownstreamStackBusLane[48][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane5_strm1_data_valid    ( DownstreamStackBusLane[48][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane6_strm0_ready         ( DownstreamStackBusLane[48][6].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane6_strm0_cntl          ( DownstreamStackBusLane[48][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane6_strm0_data          ( DownstreamStackBusLane[48][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane6_strm0_data_valid    ( DownstreamStackBusLane[48][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane6_strm1_ready         ( DownstreamStackBusLane[48][6].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane6_strm1_cntl          ( DownstreamStackBusLane[48][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane6_strm1_data          ( DownstreamStackBusLane[48][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane6_strm1_data_valid    ( DownstreamStackBusLane[48][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane7_strm0_ready         ( DownstreamStackBusLane[48][7].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane7_strm0_cntl          ( DownstreamStackBusLane[48][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane7_strm0_data          ( DownstreamStackBusLane[48][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane7_strm0_data_valid    ( DownstreamStackBusLane[48][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane7_strm1_ready         ( DownstreamStackBusLane[48][7].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane7_strm1_cntl          ( DownstreamStackBusLane[48][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane7_strm1_data          ( DownstreamStackBusLane[48][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane7_strm1_data_valid    ( DownstreamStackBusLane[48][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane8_strm0_ready         ( DownstreamStackBusLane[48][8].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane8_strm0_cntl          ( DownstreamStackBusLane[48][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane8_strm0_data          ( DownstreamStackBusLane[48][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane8_strm0_data_valid    ( DownstreamStackBusLane[48][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane8_strm1_ready         ( DownstreamStackBusLane[48][8].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane8_strm1_cntl          ( DownstreamStackBusLane[48][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane8_strm1_data          ( DownstreamStackBusLane[48][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane8_strm1_data_valid    ( DownstreamStackBusLane[48][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane9_strm0_ready         ( DownstreamStackBusLane[48][9].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane9_strm0_cntl          ( DownstreamStackBusLane[48][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane9_strm0_data          ( DownstreamStackBusLane[48][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane9_strm0_data_valid    ( DownstreamStackBusLane[48][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane9_strm1_ready         ( DownstreamStackBusLane[48][9].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane9_strm1_cntl          ( DownstreamStackBusLane[48][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane9_strm1_data          ( DownstreamStackBusLane[48][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane9_strm1_data_valid    ( DownstreamStackBusLane[48][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane10_strm0_ready         ( DownstreamStackBusLane[48][10].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane10_strm0_cntl          ( DownstreamStackBusLane[48][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane10_strm0_data          ( DownstreamStackBusLane[48][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane10_strm0_data_valid    ( DownstreamStackBusLane[48][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane10_strm1_ready         ( DownstreamStackBusLane[48][10].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane10_strm1_cntl          ( DownstreamStackBusLane[48][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane10_strm1_data          ( DownstreamStackBusLane[48][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane10_strm1_data_valid    ( DownstreamStackBusLane[48][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane11_strm0_ready         ( DownstreamStackBusLane[48][11].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane11_strm0_cntl          ( DownstreamStackBusLane[48][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane11_strm0_data          ( DownstreamStackBusLane[48][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane11_strm0_data_valid    ( DownstreamStackBusLane[48][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane11_strm1_ready         ( DownstreamStackBusLane[48][11].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane11_strm1_cntl          ( DownstreamStackBusLane[48][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane11_strm1_data          ( DownstreamStackBusLane[48][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane11_strm1_data_valid    ( DownstreamStackBusLane[48][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane12_strm0_ready         ( DownstreamStackBusLane[48][12].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane12_strm0_cntl          ( DownstreamStackBusLane[48][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane12_strm0_data          ( DownstreamStackBusLane[48][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane12_strm0_data_valid    ( DownstreamStackBusLane[48][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane12_strm1_ready         ( DownstreamStackBusLane[48][12].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane12_strm1_cntl          ( DownstreamStackBusLane[48][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane12_strm1_data          ( DownstreamStackBusLane[48][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane12_strm1_data_valid    ( DownstreamStackBusLane[48][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane13_strm0_ready         ( DownstreamStackBusLane[48][13].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane13_strm0_cntl          ( DownstreamStackBusLane[48][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane13_strm0_data          ( DownstreamStackBusLane[48][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane13_strm0_data_valid    ( DownstreamStackBusLane[48][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane13_strm1_ready         ( DownstreamStackBusLane[48][13].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane13_strm1_cntl          ( DownstreamStackBusLane[48][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane13_strm1_data          ( DownstreamStackBusLane[48][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane13_strm1_data_valid    ( DownstreamStackBusLane[48][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane14_strm0_ready         ( DownstreamStackBusLane[48][14].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane14_strm0_cntl          ( DownstreamStackBusLane[48][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane14_strm0_data          ( DownstreamStackBusLane[48][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane14_strm0_data_valid    ( DownstreamStackBusLane[48][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane14_strm1_ready         ( DownstreamStackBusLane[48][14].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane14_strm1_cntl          ( DownstreamStackBusLane[48][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane14_strm1_data          ( DownstreamStackBusLane[48][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane14_strm1_data_valid    ( DownstreamStackBusLane[48][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane15_strm0_ready         ( DownstreamStackBusLane[48][15].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane15_strm0_cntl          ( DownstreamStackBusLane[48][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane15_strm0_data          ( DownstreamStackBusLane[48][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane15_strm0_data_valid    ( DownstreamStackBusLane[48][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane15_strm1_ready         ( DownstreamStackBusLane[48][15].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane15_strm1_cntl          ( DownstreamStackBusLane[48][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane15_strm1_data          ( DownstreamStackBusLane[48][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane15_strm1_data_valid    ( DownstreamStackBusLane[48][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane16_strm0_ready         ( DownstreamStackBusLane[48][16].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane16_strm0_cntl          ( DownstreamStackBusLane[48][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane16_strm0_data          ( DownstreamStackBusLane[48][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane16_strm0_data_valid    ( DownstreamStackBusLane[48][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane16_strm1_ready         ( DownstreamStackBusLane[48][16].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane16_strm1_cntl          ( DownstreamStackBusLane[48][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane16_strm1_data          ( DownstreamStackBusLane[48][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane16_strm1_data_valid    ( DownstreamStackBusLane[48][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane17_strm0_ready         ( DownstreamStackBusLane[48][17].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane17_strm0_cntl          ( DownstreamStackBusLane[48][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane17_strm0_data          ( DownstreamStackBusLane[48][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane17_strm0_data_valid    ( DownstreamStackBusLane[48][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane17_strm1_ready         ( DownstreamStackBusLane[48][17].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane17_strm1_cntl          ( DownstreamStackBusLane[48][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane17_strm1_data          ( DownstreamStackBusLane[48][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane17_strm1_data_valid    ( DownstreamStackBusLane[48][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane18_strm0_ready         ( DownstreamStackBusLane[48][18].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane18_strm0_cntl          ( DownstreamStackBusLane[48][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane18_strm0_data          ( DownstreamStackBusLane[48][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane18_strm0_data_valid    ( DownstreamStackBusLane[48][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane18_strm1_ready         ( DownstreamStackBusLane[48][18].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane18_strm1_cntl          ( DownstreamStackBusLane[48][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane18_strm1_data          ( DownstreamStackBusLane[48][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane18_strm1_data_valid    ( DownstreamStackBusLane[48][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane19_strm0_ready         ( DownstreamStackBusLane[48][19].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane19_strm0_cntl          ( DownstreamStackBusLane[48][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane19_strm0_data          ( DownstreamStackBusLane[48][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane19_strm0_data_valid    ( DownstreamStackBusLane[48][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane19_strm1_ready         ( DownstreamStackBusLane[48][19].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane19_strm1_cntl          ( DownstreamStackBusLane[48][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane19_strm1_data          ( DownstreamStackBusLane[48][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane19_strm1_data_valid    ( DownstreamStackBusLane[48][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane20_strm0_ready         ( DownstreamStackBusLane[48][20].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane20_strm0_cntl          ( DownstreamStackBusLane[48][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane20_strm0_data          ( DownstreamStackBusLane[48][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane20_strm0_data_valid    ( DownstreamStackBusLane[48][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane20_strm1_ready         ( DownstreamStackBusLane[48][20].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane20_strm1_cntl          ( DownstreamStackBusLane[48][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane20_strm1_data          ( DownstreamStackBusLane[48][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane20_strm1_data_valid    ( DownstreamStackBusLane[48][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane21_strm0_ready         ( DownstreamStackBusLane[48][21].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane21_strm0_cntl          ( DownstreamStackBusLane[48][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane21_strm0_data          ( DownstreamStackBusLane[48][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane21_strm0_data_valid    ( DownstreamStackBusLane[48][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane21_strm1_ready         ( DownstreamStackBusLane[48][21].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane21_strm1_cntl          ( DownstreamStackBusLane[48][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane21_strm1_data          ( DownstreamStackBusLane[48][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane21_strm1_data_valid    ( DownstreamStackBusLane[48][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane22_strm0_ready         ( DownstreamStackBusLane[48][22].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane22_strm0_cntl          ( DownstreamStackBusLane[48][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane22_strm0_data          ( DownstreamStackBusLane[48][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane22_strm0_data_valid    ( DownstreamStackBusLane[48][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane22_strm1_ready         ( DownstreamStackBusLane[48][22].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane22_strm1_cntl          ( DownstreamStackBusLane[48][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane22_strm1_data          ( DownstreamStackBusLane[48][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane22_strm1_data_valid    ( DownstreamStackBusLane[48][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane23_strm0_ready         ( DownstreamStackBusLane[48][23].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane23_strm0_cntl          ( DownstreamStackBusLane[48][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane23_strm0_data          ( DownstreamStackBusLane[48][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane23_strm0_data_valid    ( DownstreamStackBusLane[48][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane23_strm1_ready         ( DownstreamStackBusLane[48][23].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane23_strm1_cntl          ( DownstreamStackBusLane[48][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane23_strm1_data          ( DownstreamStackBusLane[48][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane23_strm1_data_valid    ( DownstreamStackBusLane[48][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane24_strm0_ready         ( DownstreamStackBusLane[48][24].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane24_strm0_cntl          ( DownstreamStackBusLane[48][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane24_strm0_data          ( DownstreamStackBusLane[48][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane24_strm0_data_valid    ( DownstreamStackBusLane[48][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane24_strm1_ready         ( DownstreamStackBusLane[48][24].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane24_strm1_cntl          ( DownstreamStackBusLane[48][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane24_strm1_data          ( DownstreamStackBusLane[48][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane24_strm1_data_valid    ( DownstreamStackBusLane[48][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane25_strm0_ready         ( DownstreamStackBusLane[48][25].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane25_strm0_cntl          ( DownstreamStackBusLane[48][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane25_strm0_data          ( DownstreamStackBusLane[48][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane25_strm0_data_valid    ( DownstreamStackBusLane[48][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane25_strm1_ready         ( DownstreamStackBusLane[48][25].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane25_strm1_cntl          ( DownstreamStackBusLane[48][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane25_strm1_data          ( DownstreamStackBusLane[48][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane25_strm1_data_valid    ( DownstreamStackBusLane[48][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane26_strm0_ready         ( DownstreamStackBusLane[48][26].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane26_strm0_cntl          ( DownstreamStackBusLane[48][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane26_strm0_data          ( DownstreamStackBusLane[48][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane26_strm0_data_valid    ( DownstreamStackBusLane[48][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane26_strm1_ready         ( DownstreamStackBusLane[48][26].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane26_strm1_cntl          ( DownstreamStackBusLane[48][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane26_strm1_data          ( DownstreamStackBusLane[48][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane26_strm1_data_valid    ( DownstreamStackBusLane[48][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane27_strm0_ready         ( DownstreamStackBusLane[48][27].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane27_strm0_cntl          ( DownstreamStackBusLane[48][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane27_strm0_data          ( DownstreamStackBusLane[48][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane27_strm0_data_valid    ( DownstreamStackBusLane[48][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane27_strm1_ready         ( DownstreamStackBusLane[48][27].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane27_strm1_cntl          ( DownstreamStackBusLane[48][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane27_strm1_data          ( DownstreamStackBusLane[48][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane27_strm1_data_valid    ( DownstreamStackBusLane[48][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane28_strm0_ready         ( DownstreamStackBusLane[48][28].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane28_strm0_cntl          ( DownstreamStackBusLane[48][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane28_strm0_data          ( DownstreamStackBusLane[48][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane28_strm0_data_valid    ( DownstreamStackBusLane[48][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane28_strm1_ready         ( DownstreamStackBusLane[48][28].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane28_strm1_cntl          ( DownstreamStackBusLane[48][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane28_strm1_data          ( DownstreamStackBusLane[48][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane28_strm1_data_valid    ( DownstreamStackBusLane[48][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane29_strm0_ready         ( DownstreamStackBusLane[48][29].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane29_strm0_cntl          ( DownstreamStackBusLane[48][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane29_strm0_data          ( DownstreamStackBusLane[48][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane29_strm0_data_valid    ( DownstreamStackBusLane[48][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane29_strm1_ready         ( DownstreamStackBusLane[48][29].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane29_strm1_cntl          ( DownstreamStackBusLane[48][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane29_strm1_data          ( DownstreamStackBusLane[48][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane29_strm1_data_valid    ( DownstreamStackBusLane[48][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane30_strm0_ready         ( DownstreamStackBusLane[48][30].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane30_strm0_cntl          ( DownstreamStackBusLane[48][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane30_strm0_data          ( DownstreamStackBusLane[48][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane30_strm0_data_valid    ( DownstreamStackBusLane[48][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane30_strm1_ready         ( DownstreamStackBusLane[48][30].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane30_strm1_cntl          ( DownstreamStackBusLane[48][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane30_strm1_data          ( DownstreamStackBusLane[48][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane30_strm1_data_valid    ( DownstreamStackBusLane[48][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 48, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane31_strm0_ready         ( DownstreamStackBusLane[48][31].pe__std__lane_strm0_ready              ),      
        .std__pe48__lane31_strm0_cntl          ( DownstreamStackBusLane[48][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe48__lane31_strm0_data          ( DownstreamStackBusLane[48][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe48__lane31_strm0_data_valid    ( DownstreamStackBusLane[48][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__std__lane31_strm1_ready         ( DownstreamStackBusLane[48][31].pe__std__lane_strm1_ready              ),      
        .std__pe48__lane31_strm1_cntl          ( DownstreamStackBusLane[48][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe48__lane31_strm1_data          ( DownstreamStackBusLane[48][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe48__lane31_strm1_data_valid    ( DownstreamStackBusLane[48][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane0_strm0_ready         ( DownstreamStackBusLane[49][0].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane0_strm0_cntl          ( DownstreamStackBusLane[49][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane0_strm0_data          ( DownstreamStackBusLane[49][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane0_strm0_data_valid    ( DownstreamStackBusLane[49][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane0_strm1_ready         ( DownstreamStackBusLane[49][0].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane0_strm1_cntl          ( DownstreamStackBusLane[49][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane0_strm1_data          ( DownstreamStackBusLane[49][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane0_strm1_data_valid    ( DownstreamStackBusLane[49][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane1_strm0_ready         ( DownstreamStackBusLane[49][1].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane1_strm0_cntl          ( DownstreamStackBusLane[49][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane1_strm0_data          ( DownstreamStackBusLane[49][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane1_strm0_data_valid    ( DownstreamStackBusLane[49][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane1_strm1_ready         ( DownstreamStackBusLane[49][1].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane1_strm1_cntl          ( DownstreamStackBusLane[49][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane1_strm1_data          ( DownstreamStackBusLane[49][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane1_strm1_data_valid    ( DownstreamStackBusLane[49][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane2_strm0_ready         ( DownstreamStackBusLane[49][2].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane2_strm0_cntl          ( DownstreamStackBusLane[49][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane2_strm0_data          ( DownstreamStackBusLane[49][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane2_strm0_data_valid    ( DownstreamStackBusLane[49][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane2_strm1_ready         ( DownstreamStackBusLane[49][2].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane2_strm1_cntl          ( DownstreamStackBusLane[49][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane2_strm1_data          ( DownstreamStackBusLane[49][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane2_strm1_data_valid    ( DownstreamStackBusLane[49][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane3_strm0_ready         ( DownstreamStackBusLane[49][3].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane3_strm0_cntl          ( DownstreamStackBusLane[49][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane3_strm0_data          ( DownstreamStackBusLane[49][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane3_strm0_data_valid    ( DownstreamStackBusLane[49][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane3_strm1_ready         ( DownstreamStackBusLane[49][3].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane3_strm1_cntl          ( DownstreamStackBusLane[49][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane3_strm1_data          ( DownstreamStackBusLane[49][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane3_strm1_data_valid    ( DownstreamStackBusLane[49][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane4_strm0_ready         ( DownstreamStackBusLane[49][4].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane4_strm0_cntl          ( DownstreamStackBusLane[49][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane4_strm0_data          ( DownstreamStackBusLane[49][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane4_strm0_data_valid    ( DownstreamStackBusLane[49][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane4_strm1_ready         ( DownstreamStackBusLane[49][4].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane4_strm1_cntl          ( DownstreamStackBusLane[49][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane4_strm1_data          ( DownstreamStackBusLane[49][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane4_strm1_data_valid    ( DownstreamStackBusLane[49][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane5_strm0_ready         ( DownstreamStackBusLane[49][5].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane5_strm0_cntl          ( DownstreamStackBusLane[49][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane5_strm0_data          ( DownstreamStackBusLane[49][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane5_strm0_data_valid    ( DownstreamStackBusLane[49][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane5_strm1_ready         ( DownstreamStackBusLane[49][5].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane5_strm1_cntl          ( DownstreamStackBusLane[49][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane5_strm1_data          ( DownstreamStackBusLane[49][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane5_strm1_data_valid    ( DownstreamStackBusLane[49][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane6_strm0_ready         ( DownstreamStackBusLane[49][6].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane6_strm0_cntl          ( DownstreamStackBusLane[49][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane6_strm0_data          ( DownstreamStackBusLane[49][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane6_strm0_data_valid    ( DownstreamStackBusLane[49][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane6_strm1_ready         ( DownstreamStackBusLane[49][6].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane6_strm1_cntl          ( DownstreamStackBusLane[49][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane6_strm1_data          ( DownstreamStackBusLane[49][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane6_strm1_data_valid    ( DownstreamStackBusLane[49][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane7_strm0_ready         ( DownstreamStackBusLane[49][7].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane7_strm0_cntl          ( DownstreamStackBusLane[49][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane7_strm0_data          ( DownstreamStackBusLane[49][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane7_strm0_data_valid    ( DownstreamStackBusLane[49][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane7_strm1_ready         ( DownstreamStackBusLane[49][7].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane7_strm1_cntl          ( DownstreamStackBusLane[49][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane7_strm1_data          ( DownstreamStackBusLane[49][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane7_strm1_data_valid    ( DownstreamStackBusLane[49][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane8_strm0_ready         ( DownstreamStackBusLane[49][8].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane8_strm0_cntl          ( DownstreamStackBusLane[49][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane8_strm0_data          ( DownstreamStackBusLane[49][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane8_strm0_data_valid    ( DownstreamStackBusLane[49][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane8_strm1_ready         ( DownstreamStackBusLane[49][8].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane8_strm1_cntl          ( DownstreamStackBusLane[49][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane8_strm1_data          ( DownstreamStackBusLane[49][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane8_strm1_data_valid    ( DownstreamStackBusLane[49][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane9_strm0_ready         ( DownstreamStackBusLane[49][9].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane9_strm0_cntl          ( DownstreamStackBusLane[49][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane9_strm0_data          ( DownstreamStackBusLane[49][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane9_strm0_data_valid    ( DownstreamStackBusLane[49][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane9_strm1_ready         ( DownstreamStackBusLane[49][9].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane9_strm1_cntl          ( DownstreamStackBusLane[49][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane9_strm1_data          ( DownstreamStackBusLane[49][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane9_strm1_data_valid    ( DownstreamStackBusLane[49][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane10_strm0_ready         ( DownstreamStackBusLane[49][10].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane10_strm0_cntl          ( DownstreamStackBusLane[49][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane10_strm0_data          ( DownstreamStackBusLane[49][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane10_strm0_data_valid    ( DownstreamStackBusLane[49][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane10_strm1_ready         ( DownstreamStackBusLane[49][10].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane10_strm1_cntl          ( DownstreamStackBusLane[49][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane10_strm1_data          ( DownstreamStackBusLane[49][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane10_strm1_data_valid    ( DownstreamStackBusLane[49][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane11_strm0_ready         ( DownstreamStackBusLane[49][11].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane11_strm0_cntl          ( DownstreamStackBusLane[49][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane11_strm0_data          ( DownstreamStackBusLane[49][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane11_strm0_data_valid    ( DownstreamStackBusLane[49][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane11_strm1_ready         ( DownstreamStackBusLane[49][11].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane11_strm1_cntl          ( DownstreamStackBusLane[49][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane11_strm1_data          ( DownstreamStackBusLane[49][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane11_strm1_data_valid    ( DownstreamStackBusLane[49][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane12_strm0_ready         ( DownstreamStackBusLane[49][12].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane12_strm0_cntl          ( DownstreamStackBusLane[49][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane12_strm0_data          ( DownstreamStackBusLane[49][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane12_strm0_data_valid    ( DownstreamStackBusLane[49][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane12_strm1_ready         ( DownstreamStackBusLane[49][12].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane12_strm1_cntl          ( DownstreamStackBusLane[49][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane12_strm1_data          ( DownstreamStackBusLane[49][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane12_strm1_data_valid    ( DownstreamStackBusLane[49][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane13_strm0_ready         ( DownstreamStackBusLane[49][13].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane13_strm0_cntl          ( DownstreamStackBusLane[49][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane13_strm0_data          ( DownstreamStackBusLane[49][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane13_strm0_data_valid    ( DownstreamStackBusLane[49][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane13_strm1_ready         ( DownstreamStackBusLane[49][13].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane13_strm1_cntl          ( DownstreamStackBusLane[49][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane13_strm1_data          ( DownstreamStackBusLane[49][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane13_strm1_data_valid    ( DownstreamStackBusLane[49][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane14_strm0_ready         ( DownstreamStackBusLane[49][14].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane14_strm0_cntl          ( DownstreamStackBusLane[49][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane14_strm0_data          ( DownstreamStackBusLane[49][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane14_strm0_data_valid    ( DownstreamStackBusLane[49][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane14_strm1_ready         ( DownstreamStackBusLane[49][14].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane14_strm1_cntl          ( DownstreamStackBusLane[49][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane14_strm1_data          ( DownstreamStackBusLane[49][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane14_strm1_data_valid    ( DownstreamStackBusLane[49][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane15_strm0_ready         ( DownstreamStackBusLane[49][15].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane15_strm0_cntl          ( DownstreamStackBusLane[49][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane15_strm0_data          ( DownstreamStackBusLane[49][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane15_strm0_data_valid    ( DownstreamStackBusLane[49][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane15_strm1_ready         ( DownstreamStackBusLane[49][15].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane15_strm1_cntl          ( DownstreamStackBusLane[49][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane15_strm1_data          ( DownstreamStackBusLane[49][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane15_strm1_data_valid    ( DownstreamStackBusLane[49][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane16_strm0_ready         ( DownstreamStackBusLane[49][16].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane16_strm0_cntl          ( DownstreamStackBusLane[49][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane16_strm0_data          ( DownstreamStackBusLane[49][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane16_strm0_data_valid    ( DownstreamStackBusLane[49][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane16_strm1_ready         ( DownstreamStackBusLane[49][16].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane16_strm1_cntl          ( DownstreamStackBusLane[49][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane16_strm1_data          ( DownstreamStackBusLane[49][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane16_strm1_data_valid    ( DownstreamStackBusLane[49][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane17_strm0_ready         ( DownstreamStackBusLane[49][17].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane17_strm0_cntl          ( DownstreamStackBusLane[49][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane17_strm0_data          ( DownstreamStackBusLane[49][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane17_strm0_data_valid    ( DownstreamStackBusLane[49][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane17_strm1_ready         ( DownstreamStackBusLane[49][17].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane17_strm1_cntl          ( DownstreamStackBusLane[49][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane17_strm1_data          ( DownstreamStackBusLane[49][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane17_strm1_data_valid    ( DownstreamStackBusLane[49][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane18_strm0_ready         ( DownstreamStackBusLane[49][18].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane18_strm0_cntl          ( DownstreamStackBusLane[49][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane18_strm0_data          ( DownstreamStackBusLane[49][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane18_strm0_data_valid    ( DownstreamStackBusLane[49][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane18_strm1_ready         ( DownstreamStackBusLane[49][18].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane18_strm1_cntl          ( DownstreamStackBusLane[49][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane18_strm1_data          ( DownstreamStackBusLane[49][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane18_strm1_data_valid    ( DownstreamStackBusLane[49][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane19_strm0_ready         ( DownstreamStackBusLane[49][19].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane19_strm0_cntl          ( DownstreamStackBusLane[49][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane19_strm0_data          ( DownstreamStackBusLane[49][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane19_strm0_data_valid    ( DownstreamStackBusLane[49][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane19_strm1_ready         ( DownstreamStackBusLane[49][19].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane19_strm1_cntl          ( DownstreamStackBusLane[49][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane19_strm1_data          ( DownstreamStackBusLane[49][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane19_strm1_data_valid    ( DownstreamStackBusLane[49][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane20_strm0_ready         ( DownstreamStackBusLane[49][20].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane20_strm0_cntl          ( DownstreamStackBusLane[49][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane20_strm0_data          ( DownstreamStackBusLane[49][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane20_strm0_data_valid    ( DownstreamStackBusLane[49][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane20_strm1_ready         ( DownstreamStackBusLane[49][20].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane20_strm1_cntl          ( DownstreamStackBusLane[49][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane20_strm1_data          ( DownstreamStackBusLane[49][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane20_strm1_data_valid    ( DownstreamStackBusLane[49][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane21_strm0_ready         ( DownstreamStackBusLane[49][21].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane21_strm0_cntl          ( DownstreamStackBusLane[49][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane21_strm0_data          ( DownstreamStackBusLane[49][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane21_strm0_data_valid    ( DownstreamStackBusLane[49][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane21_strm1_ready         ( DownstreamStackBusLane[49][21].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane21_strm1_cntl          ( DownstreamStackBusLane[49][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane21_strm1_data          ( DownstreamStackBusLane[49][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane21_strm1_data_valid    ( DownstreamStackBusLane[49][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane22_strm0_ready         ( DownstreamStackBusLane[49][22].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane22_strm0_cntl          ( DownstreamStackBusLane[49][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane22_strm0_data          ( DownstreamStackBusLane[49][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane22_strm0_data_valid    ( DownstreamStackBusLane[49][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane22_strm1_ready         ( DownstreamStackBusLane[49][22].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane22_strm1_cntl          ( DownstreamStackBusLane[49][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane22_strm1_data          ( DownstreamStackBusLane[49][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane22_strm1_data_valid    ( DownstreamStackBusLane[49][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane23_strm0_ready         ( DownstreamStackBusLane[49][23].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane23_strm0_cntl          ( DownstreamStackBusLane[49][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane23_strm0_data          ( DownstreamStackBusLane[49][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane23_strm0_data_valid    ( DownstreamStackBusLane[49][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane23_strm1_ready         ( DownstreamStackBusLane[49][23].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane23_strm1_cntl          ( DownstreamStackBusLane[49][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane23_strm1_data          ( DownstreamStackBusLane[49][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane23_strm1_data_valid    ( DownstreamStackBusLane[49][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane24_strm0_ready         ( DownstreamStackBusLane[49][24].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane24_strm0_cntl          ( DownstreamStackBusLane[49][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane24_strm0_data          ( DownstreamStackBusLane[49][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane24_strm0_data_valid    ( DownstreamStackBusLane[49][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane24_strm1_ready         ( DownstreamStackBusLane[49][24].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane24_strm1_cntl          ( DownstreamStackBusLane[49][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane24_strm1_data          ( DownstreamStackBusLane[49][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane24_strm1_data_valid    ( DownstreamStackBusLane[49][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane25_strm0_ready         ( DownstreamStackBusLane[49][25].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane25_strm0_cntl          ( DownstreamStackBusLane[49][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane25_strm0_data          ( DownstreamStackBusLane[49][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane25_strm0_data_valid    ( DownstreamStackBusLane[49][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane25_strm1_ready         ( DownstreamStackBusLane[49][25].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane25_strm1_cntl          ( DownstreamStackBusLane[49][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane25_strm1_data          ( DownstreamStackBusLane[49][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane25_strm1_data_valid    ( DownstreamStackBusLane[49][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane26_strm0_ready         ( DownstreamStackBusLane[49][26].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane26_strm0_cntl          ( DownstreamStackBusLane[49][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane26_strm0_data          ( DownstreamStackBusLane[49][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane26_strm0_data_valid    ( DownstreamStackBusLane[49][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane26_strm1_ready         ( DownstreamStackBusLane[49][26].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane26_strm1_cntl          ( DownstreamStackBusLane[49][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane26_strm1_data          ( DownstreamStackBusLane[49][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane26_strm1_data_valid    ( DownstreamStackBusLane[49][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane27_strm0_ready         ( DownstreamStackBusLane[49][27].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane27_strm0_cntl          ( DownstreamStackBusLane[49][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane27_strm0_data          ( DownstreamStackBusLane[49][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane27_strm0_data_valid    ( DownstreamStackBusLane[49][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane27_strm1_ready         ( DownstreamStackBusLane[49][27].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane27_strm1_cntl          ( DownstreamStackBusLane[49][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane27_strm1_data          ( DownstreamStackBusLane[49][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane27_strm1_data_valid    ( DownstreamStackBusLane[49][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane28_strm0_ready         ( DownstreamStackBusLane[49][28].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane28_strm0_cntl          ( DownstreamStackBusLane[49][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane28_strm0_data          ( DownstreamStackBusLane[49][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane28_strm0_data_valid    ( DownstreamStackBusLane[49][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane28_strm1_ready         ( DownstreamStackBusLane[49][28].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane28_strm1_cntl          ( DownstreamStackBusLane[49][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane28_strm1_data          ( DownstreamStackBusLane[49][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane28_strm1_data_valid    ( DownstreamStackBusLane[49][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane29_strm0_ready         ( DownstreamStackBusLane[49][29].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane29_strm0_cntl          ( DownstreamStackBusLane[49][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane29_strm0_data          ( DownstreamStackBusLane[49][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane29_strm0_data_valid    ( DownstreamStackBusLane[49][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane29_strm1_ready         ( DownstreamStackBusLane[49][29].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane29_strm1_cntl          ( DownstreamStackBusLane[49][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane29_strm1_data          ( DownstreamStackBusLane[49][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane29_strm1_data_valid    ( DownstreamStackBusLane[49][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane30_strm0_ready         ( DownstreamStackBusLane[49][30].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane30_strm0_cntl          ( DownstreamStackBusLane[49][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane30_strm0_data          ( DownstreamStackBusLane[49][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane30_strm0_data_valid    ( DownstreamStackBusLane[49][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane30_strm1_ready         ( DownstreamStackBusLane[49][30].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane30_strm1_cntl          ( DownstreamStackBusLane[49][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane30_strm1_data          ( DownstreamStackBusLane[49][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane30_strm1_data_valid    ( DownstreamStackBusLane[49][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 49, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane31_strm0_ready         ( DownstreamStackBusLane[49][31].pe__std__lane_strm0_ready              ),      
        .std__pe49__lane31_strm0_cntl          ( DownstreamStackBusLane[49][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe49__lane31_strm0_data          ( DownstreamStackBusLane[49][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe49__lane31_strm0_data_valid    ( DownstreamStackBusLane[49][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__std__lane31_strm1_ready         ( DownstreamStackBusLane[49][31].pe__std__lane_strm1_ready              ),      
        .std__pe49__lane31_strm1_cntl          ( DownstreamStackBusLane[49][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe49__lane31_strm1_data          ( DownstreamStackBusLane[49][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe49__lane31_strm1_data_valid    ( DownstreamStackBusLane[49][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane0_strm0_ready         ( DownstreamStackBusLane[50][0].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane0_strm0_cntl          ( DownstreamStackBusLane[50][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane0_strm0_data          ( DownstreamStackBusLane[50][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane0_strm0_data_valid    ( DownstreamStackBusLane[50][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane0_strm1_ready         ( DownstreamStackBusLane[50][0].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane0_strm1_cntl          ( DownstreamStackBusLane[50][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane0_strm1_data          ( DownstreamStackBusLane[50][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane0_strm1_data_valid    ( DownstreamStackBusLane[50][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane1_strm0_ready         ( DownstreamStackBusLane[50][1].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane1_strm0_cntl          ( DownstreamStackBusLane[50][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane1_strm0_data          ( DownstreamStackBusLane[50][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane1_strm0_data_valid    ( DownstreamStackBusLane[50][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane1_strm1_ready         ( DownstreamStackBusLane[50][1].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane1_strm1_cntl          ( DownstreamStackBusLane[50][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane1_strm1_data          ( DownstreamStackBusLane[50][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane1_strm1_data_valid    ( DownstreamStackBusLane[50][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane2_strm0_ready         ( DownstreamStackBusLane[50][2].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane2_strm0_cntl          ( DownstreamStackBusLane[50][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane2_strm0_data          ( DownstreamStackBusLane[50][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane2_strm0_data_valid    ( DownstreamStackBusLane[50][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane2_strm1_ready         ( DownstreamStackBusLane[50][2].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane2_strm1_cntl          ( DownstreamStackBusLane[50][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane2_strm1_data          ( DownstreamStackBusLane[50][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane2_strm1_data_valid    ( DownstreamStackBusLane[50][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane3_strm0_ready         ( DownstreamStackBusLane[50][3].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane3_strm0_cntl          ( DownstreamStackBusLane[50][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane3_strm0_data          ( DownstreamStackBusLane[50][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane3_strm0_data_valid    ( DownstreamStackBusLane[50][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane3_strm1_ready         ( DownstreamStackBusLane[50][3].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane3_strm1_cntl          ( DownstreamStackBusLane[50][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane3_strm1_data          ( DownstreamStackBusLane[50][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane3_strm1_data_valid    ( DownstreamStackBusLane[50][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane4_strm0_ready         ( DownstreamStackBusLane[50][4].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane4_strm0_cntl          ( DownstreamStackBusLane[50][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane4_strm0_data          ( DownstreamStackBusLane[50][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane4_strm0_data_valid    ( DownstreamStackBusLane[50][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane4_strm1_ready         ( DownstreamStackBusLane[50][4].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane4_strm1_cntl          ( DownstreamStackBusLane[50][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane4_strm1_data          ( DownstreamStackBusLane[50][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane4_strm1_data_valid    ( DownstreamStackBusLane[50][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane5_strm0_ready         ( DownstreamStackBusLane[50][5].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane5_strm0_cntl          ( DownstreamStackBusLane[50][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane5_strm0_data          ( DownstreamStackBusLane[50][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane5_strm0_data_valid    ( DownstreamStackBusLane[50][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane5_strm1_ready         ( DownstreamStackBusLane[50][5].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane5_strm1_cntl          ( DownstreamStackBusLane[50][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane5_strm1_data          ( DownstreamStackBusLane[50][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane5_strm1_data_valid    ( DownstreamStackBusLane[50][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane6_strm0_ready         ( DownstreamStackBusLane[50][6].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane6_strm0_cntl          ( DownstreamStackBusLane[50][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane6_strm0_data          ( DownstreamStackBusLane[50][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane6_strm0_data_valid    ( DownstreamStackBusLane[50][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane6_strm1_ready         ( DownstreamStackBusLane[50][6].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane6_strm1_cntl          ( DownstreamStackBusLane[50][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane6_strm1_data          ( DownstreamStackBusLane[50][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane6_strm1_data_valid    ( DownstreamStackBusLane[50][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane7_strm0_ready         ( DownstreamStackBusLane[50][7].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane7_strm0_cntl          ( DownstreamStackBusLane[50][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane7_strm0_data          ( DownstreamStackBusLane[50][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane7_strm0_data_valid    ( DownstreamStackBusLane[50][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane7_strm1_ready         ( DownstreamStackBusLane[50][7].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane7_strm1_cntl          ( DownstreamStackBusLane[50][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane7_strm1_data          ( DownstreamStackBusLane[50][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane7_strm1_data_valid    ( DownstreamStackBusLane[50][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane8_strm0_ready         ( DownstreamStackBusLane[50][8].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane8_strm0_cntl          ( DownstreamStackBusLane[50][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane8_strm0_data          ( DownstreamStackBusLane[50][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane8_strm0_data_valid    ( DownstreamStackBusLane[50][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane8_strm1_ready         ( DownstreamStackBusLane[50][8].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane8_strm1_cntl          ( DownstreamStackBusLane[50][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane8_strm1_data          ( DownstreamStackBusLane[50][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane8_strm1_data_valid    ( DownstreamStackBusLane[50][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane9_strm0_ready         ( DownstreamStackBusLane[50][9].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane9_strm0_cntl          ( DownstreamStackBusLane[50][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane9_strm0_data          ( DownstreamStackBusLane[50][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane9_strm0_data_valid    ( DownstreamStackBusLane[50][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane9_strm1_ready         ( DownstreamStackBusLane[50][9].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane9_strm1_cntl          ( DownstreamStackBusLane[50][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane9_strm1_data          ( DownstreamStackBusLane[50][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane9_strm1_data_valid    ( DownstreamStackBusLane[50][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane10_strm0_ready         ( DownstreamStackBusLane[50][10].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane10_strm0_cntl          ( DownstreamStackBusLane[50][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane10_strm0_data          ( DownstreamStackBusLane[50][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane10_strm0_data_valid    ( DownstreamStackBusLane[50][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane10_strm1_ready         ( DownstreamStackBusLane[50][10].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane10_strm1_cntl          ( DownstreamStackBusLane[50][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane10_strm1_data          ( DownstreamStackBusLane[50][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane10_strm1_data_valid    ( DownstreamStackBusLane[50][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane11_strm0_ready         ( DownstreamStackBusLane[50][11].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane11_strm0_cntl          ( DownstreamStackBusLane[50][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane11_strm0_data          ( DownstreamStackBusLane[50][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane11_strm0_data_valid    ( DownstreamStackBusLane[50][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane11_strm1_ready         ( DownstreamStackBusLane[50][11].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane11_strm1_cntl          ( DownstreamStackBusLane[50][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane11_strm1_data          ( DownstreamStackBusLane[50][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane11_strm1_data_valid    ( DownstreamStackBusLane[50][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane12_strm0_ready         ( DownstreamStackBusLane[50][12].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane12_strm0_cntl          ( DownstreamStackBusLane[50][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane12_strm0_data          ( DownstreamStackBusLane[50][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane12_strm0_data_valid    ( DownstreamStackBusLane[50][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane12_strm1_ready         ( DownstreamStackBusLane[50][12].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane12_strm1_cntl          ( DownstreamStackBusLane[50][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane12_strm1_data          ( DownstreamStackBusLane[50][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane12_strm1_data_valid    ( DownstreamStackBusLane[50][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane13_strm0_ready         ( DownstreamStackBusLane[50][13].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane13_strm0_cntl          ( DownstreamStackBusLane[50][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane13_strm0_data          ( DownstreamStackBusLane[50][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane13_strm0_data_valid    ( DownstreamStackBusLane[50][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane13_strm1_ready         ( DownstreamStackBusLane[50][13].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane13_strm1_cntl          ( DownstreamStackBusLane[50][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane13_strm1_data          ( DownstreamStackBusLane[50][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane13_strm1_data_valid    ( DownstreamStackBusLane[50][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane14_strm0_ready         ( DownstreamStackBusLane[50][14].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane14_strm0_cntl          ( DownstreamStackBusLane[50][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane14_strm0_data          ( DownstreamStackBusLane[50][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane14_strm0_data_valid    ( DownstreamStackBusLane[50][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane14_strm1_ready         ( DownstreamStackBusLane[50][14].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane14_strm1_cntl          ( DownstreamStackBusLane[50][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane14_strm1_data          ( DownstreamStackBusLane[50][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane14_strm1_data_valid    ( DownstreamStackBusLane[50][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane15_strm0_ready         ( DownstreamStackBusLane[50][15].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane15_strm0_cntl          ( DownstreamStackBusLane[50][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane15_strm0_data          ( DownstreamStackBusLane[50][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane15_strm0_data_valid    ( DownstreamStackBusLane[50][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane15_strm1_ready         ( DownstreamStackBusLane[50][15].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane15_strm1_cntl          ( DownstreamStackBusLane[50][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane15_strm1_data          ( DownstreamStackBusLane[50][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane15_strm1_data_valid    ( DownstreamStackBusLane[50][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane16_strm0_ready         ( DownstreamStackBusLane[50][16].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane16_strm0_cntl          ( DownstreamStackBusLane[50][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane16_strm0_data          ( DownstreamStackBusLane[50][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane16_strm0_data_valid    ( DownstreamStackBusLane[50][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane16_strm1_ready         ( DownstreamStackBusLane[50][16].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane16_strm1_cntl          ( DownstreamStackBusLane[50][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane16_strm1_data          ( DownstreamStackBusLane[50][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane16_strm1_data_valid    ( DownstreamStackBusLane[50][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane17_strm0_ready         ( DownstreamStackBusLane[50][17].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane17_strm0_cntl          ( DownstreamStackBusLane[50][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane17_strm0_data          ( DownstreamStackBusLane[50][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane17_strm0_data_valid    ( DownstreamStackBusLane[50][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane17_strm1_ready         ( DownstreamStackBusLane[50][17].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane17_strm1_cntl          ( DownstreamStackBusLane[50][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane17_strm1_data          ( DownstreamStackBusLane[50][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane17_strm1_data_valid    ( DownstreamStackBusLane[50][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane18_strm0_ready         ( DownstreamStackBusLane[50][18].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane18_strm0_cntl          ( DownstreamStackBusLane[50][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane18_strm0_data          ( DownstreamStackBusLane[50][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane18_strm0_data_valid    ( DownstreamStackBusLane[50][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane18_strm1_ready         ( DownstreamStackBusLane[50][18].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane18_strm1_cntl          ( DownstreamStackBusLane[50][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane18_strm1_data          ( DownstreamStackBusLane[50][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane18_strm1_data_valid    ( DownstreamStackBusLane[50][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane19_strm0_ready         ( DownstreamStackBusLane[50][19].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane19_strm0_cntl          ( DownstreamStackBusLane[50][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane19_strm0_data          ( DownstreamStackBusLane[50][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane19_strm0_data_valid    ( DownstreamStackBusLane[50][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane19_strm1_ready         ( DownstreamStackBusLane[50][19].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane19_strm1_cntl          ( DownstreamStackBusLane[50][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane19_strm1_data          ( DownstreamStackBusLane[50][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane19_strm1_data_valid    ( DownstreamStackBusLane[50][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane20_strm0_ready         ( DownstreamStackBusLane[50][20].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane20_strm0_cntl          ( DownstreamStackBusLane[50][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane20_strm0_data          ( DownstreamStackBusLane[50][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane20_strm0_data_valid    ( DownstreamStackBusLane[50][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane20_strm1_ready         ( DownstreamStackBusLane[50][20].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane20_strm1_cntl          ( DownstreamStackBusLane[50][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane20_strm1_data          ( DownstreamStackBusLane[50][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane20_strm1_data_valid    ( DownstreamStackBusLane[50][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane21_strm0_ready         ( DownstreamStackBusLane[50][21].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane21_strm0_cntl          ( DownstreamStackBusLane[50][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane21_strm0_data          ( DownstreamStackBusLane[50][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane21_strm0_data_valid    ( DownstreamStackBusLane[50][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane21_strm1_ready         ( DownstreamStackBusLane[50][21].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane21_strm1_cntl          ( DownstreamStackBusLane[50][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane21_strm1_data          ( DownstreamStackBusLane[50][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane21_strm1_data_valid    ( DownstreamStackBusLane[50][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane22_strm0_ready         ( DownstreamStackBusLane[50][22].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane22_strm0_cntl          ( DownstreamStackBusLane[50][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane22_strm0_data          ( DownstreamStackBusLane[50][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane22_strm0_data_valid    ( DownstreamStackBusLane[50][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane22_strm1_ready         ( DownstreamStackBusLane[50][22].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane22_strm1_cntl          ( DownstreamStackBusLane[50][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane22_strm1_data          ( DownstreamStackBusLane[50][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane22_strm1_data_valid    ( DownstreamStackBusLane[50][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane23_strm0_ready         ( DownstreamStackBusLane[50][23].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane23_strm0_cntl          ( DownstreamStackBusLane[50][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane23_strm0_data          ( DownstreamStackBusLane[50][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane23_strm0_data_valid    ( DownstreamStackBusLane[50][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane23_strm1_ready         ( DownstreamStackBusLane[50][23].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane23_strm1_cntl          ( DownstreamStackBusLane[50][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane23_strm1_data          ( DownstreamStackBusLane[50][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane23_strm1_data_valid    ( DownstreamStackBusLane[50][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane24_strm0_ready         ( DownstreamStackBusLane[50][24].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane24_strm0_cntl          ( DownstreamStackBusLane[50][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane24_strm0_data          ( DownstreamStackBusLane[50][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane24_strm0_data_valid    ( DownstreamStackBusLane[50][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane24_strm1_ready         ( DownstreamStackBusLane[50][24].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane24_strm1_cntl          ( DownstreamStackBusLane[50][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane24_strm1_data          ( DownstreamStackBusLane[50][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane24_strm1_data_valid    ( DownstreamStackBusLane[50][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane25_strm0_ready         ( DownstreamStackBusLane[50][25].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane25_strm0_cntl          ( DownstreamStackBusLane[50][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane25_strm0_data          ( DownstreamStackBusLane[50][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane25_strm0_data_valid    ( DownstreamStackBusLane[50][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane25_strm1_ready         ( DownstreamStackBusLane[50][25].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane25_strm1_cntl          ( DownstreamStackBusLane[50][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane25_strm1_data          ( DownstreamStackBusLane[50][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane25_strm1_data_valid    ( DownstreamStackBusLane[50][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane26_strm0_ready         ( DownstreamStackBusLane[50][26].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane26_strm0_cntl          ( DownstreamStackBusLane[50][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane26_strm0_data          ( DownstreamStackBusLane[50][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane26_strm0_data_valid    ( DownstreamStackBusLane[50][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane26_strm1_ready         ( DownstreamStackBusLane[50][26].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane26_strm1_cntl          ( DownstreamStackBusLane[50][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane26_strm1_data          ( DownstreamStackBusLane[50][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane26_strm1_data_valid    ( DownstreamStackBusLane[50][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane27_strm0_ready         ( DownstreamStackBusLane[50][27].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane27_strm0_cntl          ( DownstreamStackBusLane[50][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane27_strm0_data          ( DownstreamStackBusLane[50][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane27_strm0_data_valid    ( DownstreamStackBusLane[50][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane27_strm1_ready         ( DownstreamStackBusLane[50][27].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane27_strm1_cntl          ( DownstreamStackBusLane[50][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane27_strm1_data          ( DownstreamStackBusLane[50][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane27_strm1_data_valid    ( DownstreamStackBusLane[50][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane28_strm0_ready         ( DownstreamStackBusLane[50][28].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane28_strm0_cntl          ( DownstreamStackBusLane[50][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane28_strm0_data          ( DownstreamStackBusLane[50][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane28_strm0_data_valid    ( DownstreamStackBusLane[50][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane28_strm1_ready         ( DownstreamStackBusLane[50][28].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane28_strm1_cntl          ( DownstreamStackBusLane[50][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane28_strm1_data          ( DownstreamStackBusLane[50][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane28_strm1_data_valid    ( DownstreamStackBusLane[50][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane29_strm0_ready         ( DownstreamStackBusLane[50][29].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane29_strm0_cntl          ( DownstreamStackBusLane[50][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane29_strm0_data          ( DownstreamStackBusLane[50][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane29_strm0_data_valid    ( DownstreamStackBusLane[50][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane29_strm1_ready         ( DownstreamStackBusLane[50][29].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane29_strm1_cntl          ( DownstreamStackBusLane[50][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane29_strm1_data          ( DownstreamStackBusLane[50][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane29_strm1_data_valid    ( DownstreamStackBusLane[50][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane30_strm0_ready         ( DownstreamStackBusLane[50][30].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane30_strm0_cntl          ( DownstreamStackBusLane[50][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane30_strm0_data          ( DownstreamStackBusLane[50][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane30_strm0_data_valid    ( DownstreamStackBusLane[50][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane30_strm1_ready         ( DownstreamStackBusLane[50][30].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane30_strm1_cntl          ( DownstreamStackBusLane[50][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane30_strm1_data          ( DownstreamStackBusLane[50][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane30_strm1_data_valid    ( DownstreamStackBusLane[50][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 50, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane31_strm0_ready         ( DownstreamStackBusLane[50][31].pe__std__lane_strm0_ready              ),      
        .std__pe50__lane31_strm0_cntl          ( DownstreamStackBusLane[50][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe50__lane31_strm0_data          ( DownstreamStackBusLane[50][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe50__lane31_strm0_data_valid    ( DownstreamStackBusLane[50][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__std__lane31_strm1_ready         ( DownstreamStackBusLane[50][31].pe__std__lane_strm1_ready              ),      
        .std__pe50__lane31_strm1_cntl          ( DownstreamStackBusLane[50][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe50__lane31_strm1_data          ( DownstreamStackBusLane[50][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe50__lane31_strm1_data_valid    ( DownstreamStackBusLane[50][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane0_strm0_ready         ( DownstreamStackBusLane[51][0].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane0_strm0_cntl          ( DownstreamStackBusLane[51][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane0_strm0_data          ( DownstreamStackBusLane[51][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane0_strm0_data_valid    ( DownstreamStackBusLane[51][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane0_strm1_ready         ( DownstreamStackBusLane[51][0].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane0_strm1_cntl          ( DownstreamStackBusLane[51][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane0_strm1_data          ( DownstreamStackBusLane[51][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane0_strm1_data_valid    ( DownstreamStackBusLane[51][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane1_strm0_ready         ( DownstreamStackBusLane[51][1].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane1_strm0_cntl          ( DownstreamStackBusLane[51][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane1_strm0_data          ( DownstreamStackBusLane[51][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane1_strm0_data_valid    ( DownstreamStackBusLane[51][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane1_strm1_ready         ( DownstreamStackBusLane[51][1].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane1_strm1_cntl          ( DownstreamStackBusLane[51][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane1_strm1_data          ( DownstreamStackBusLane[51][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane1_strm1_data_valid    ( DownstreamStackBusLane[51][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane2_strm0_ready         ( DownstreamStackBusLane[51][2].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane2_strm0_cntl          ( DownstreamStackBusLane[51][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane2_strm0_data          ( DownstreamStackBusLane[51][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane2_strm0_data_valid    ( DownstreamStackBusLane[51][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane2_strm1_ready         ( DownstreamStackBusLane[51][2].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane2_strm1_cntl          ( DownstreamStackBusLane[51][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane2_strm1_data          ( DownstreamStackBusLane[51][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane2_strm1_data_valid    ( DownstreamStackBusLane[51][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane3_strm0_ready         ( DownstreamStackBusLane[51][3].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane3_strm0_cntl          ( DownstreamStackBusLane[51][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane3_strm0_data          ( DownstreamStackBusLane[51][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane3_strm0_data_valid    ( DownstreamStackBusLane[51][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane3_strm1_ready         ( DownstreamStackBusLane[51][3].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane3_strm1_cntl          ( DownstreamStackBusLane[51][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane3_strm1_data          ( DownstreamStackBusLane[51][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane3_strm1_data_valid    ( DownstreamStackBusLane[51][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane4_strm0_ready         ( DownstreamStackBusLane[51][4].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane4_strm0_cntl          ( DownstreamStackBusLane[51][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane4_strm0_data          ( DownstreamStackBusLane[51][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane4_strm0_data_valid    ( DownstreamStackBusLane[51][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane4_strm1_ready         ( DownstreamStackBusLane[51][4].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane4_strm1_cntl          ( DownstreamStackBusLane[51][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane4_strm1_data          ( DownstreamStackBusLane[51][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane4_strm1_data_valid    ( DownstreamStackBusLane[51][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane5_strm0_ready         ( DownstreamStackBusLane[51][5].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane5_strm0_cntl          ( DownstreamStackBusLane[51][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane5_strm0_data          ( DownstreamStackBusLane[51][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane5_strm0_data_valid    ( DownstreamStackBusLane[51][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane5_strm1_ready         ( DownstreamStackBusLane[51][5].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane5_strm1_cntl          ( DownstreamStackBusLane[51][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane5_strm1_data          ( DownstreamStackBusLane[51][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane5_strm1_data_valid    ( DownstreamStackBusLane[51][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane6_strm0_ready         ( DownstreamStackBusLane[51][6].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane6_strm0_cntl          ( DownstreamStackBusLane[51][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane6_strm0_data          ( DownstreamStackBusLane[51][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane6_strm0_data_valid    ( DownstreamStackBusLane[51][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane6_strm1_ready         ( DownstreamStackBusLane[51][6].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane6_strm1_cntl          ( DownstreamStackBusLane[51][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane6_strm1_data          ( DownstreamStackBusLane[51][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane6_strm1_data_valid    ( DownstreamStackBusLane[51][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane7_strm0_ready         ( DownstreamStackBusLane[51][7].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane7_strm0_cntl          ( DownstreamStackBusLane[51][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane7_strm0_data          ( DownstreamStackBusLane[51][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane7_strm0_data_valid    ( DownstreamStackBusLane[51][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane7_strm1_ready         ( DownstreamStackBusLane[51][7].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane7_strm1_cntl          ( DownstreamStackBusLane[51][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane7_strm1_data          ( DownstreamStackBusLane[51][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane7_strm1_data_valid    ( DownstreamStackBusLane[51][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane8_strm0_ready         ( DownstreamStackBusLane[51][8].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane8_strm0_cntl          ( DownstreamStackBusLane[51][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane8_strm0_data          ( DownstreamStackBusLane[51][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane8_strm0_data_valid    ( DownstreamStackBusLane[51][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane8_strm1_ready         ( DownstreamStackBusLane[51][8].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane8_strm1_cntl          ( DownstreamStackBusLane[51][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane8_strm1_data          ( DownstreamStackBusLane[51][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane8_strm1_data_valid    ( DownstreamStackBusLane[51][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane9_strm0_ready         ( DownstreamStackBusLane[51][9].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane9_strm0_cntl          ( DownstreamStackBusLane[51][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane9_strm0_data          ( DownstreamStackBusLane[51][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane9_strm0_data_valid    ( DownstreamStackBusLane[51][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane9_strm1_ready         ( DownstreamStackBusLane[51][9].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane9_strm1_cntl          ( DownstreamStackBusLane[51][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane9_strm1_data          ( DownstreamStackBusLane[51][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane9_strm1_data_valid    ( DownstreamStackBusLane[51][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane10_strm0_ready         ( DownstreamStackBusLane[51][10].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane10_strm0_cntl          ( DownstreamStackBusLane[51][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane10_strm0_data          ( DownstreamStackBusLane[51][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane10_strm0_data_valid    ( DownstreamStackBusLane[51][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane10_strm1_ready         ( DownstreamStackBusLane[51][10].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane10_strm1_cntl          ( DownstreamStackBusLane[51][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane10_strm1_data          ( DownstreamStackBusLane[51][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane10_strm1_data_valid    ( DownstreamStackBusLane[51][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane11_strm0_ready         ( DownstreamStackBusLane[51][11].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane11_strm0_cntl          ( DownstreamStackBusLane[51][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane11_strm0_data          ( DownstreamStackBusLane[51][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane11_strm0_data_valid    ( DownstreamStackBusLane[51][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane11_strm1_ready         ( DownstreamStackBusLane[51][11].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane11_strm1_cntl          ( DownstreamStackBusLane[51][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane11_strm1_data          ( DownstreamStackBusLane[51][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane11_strm1_data_valid    ( DownstreamStackBusLane[51][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane12_strm0_ready         ( DownstreamStackBusLane[51][12].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane12_strm0_cntl          ( DownstreamStackBusLane[51][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane12_strm0_data          ( DownstreamStackBusLane[51][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane12_strm0_data_valid    ( DownstreamStackBusLane[51][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane12_strm1_ready         ( DownstreamStackBusLane[51][12].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane12_strm1_cntl          ( DownstreamStackBusLane[51][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane12_strm1_data          ( DownstreamStackBusLane[51][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane12_strm1_data_valid    ( DownstreamStackBusLane[51][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane13_strm0_ready         ( DownstreamStackBusLane[51][13].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane13_strm0_cntl          ( DownstreamStackBusLane[51][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane13_strm0_data          ( DownstreamStackBusLane[51][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane13_strm0_data_valid    ( DownstreamStackBusLane[51][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane13_strm1_ready         ( DownstreamStackBusLane[51][13].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane13_strm1_cntl          ( DownstreamStackBusLane[51][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane13_strm1_data          ( DownstreamStackBusLane[51][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane13_strm1_data_valid    ( DownstreamStackBusLane[51][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane14_strm0_ready         ( DownstreamStackBusLane[51][14].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane14_strm0_cntl          ( DownstreamStackBusLane[51][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane14_strm0_data          ( DownstreamStackBusLane[51][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane14_strm0_data_valid    ( DownstreamStackBusLane[51][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane14_strm1_ready         ( DownstreamStackBusLane[51][14].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane14_strm1_cntl          ( DownstreamStackBusLane[51][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane14_strm1_data          ( DownstreamStackBusLane[51][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane14_strm1_data_valid    ( DownstreamStackBusLane[51][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane15_strm0_ready         ( DownstreamStackBusLane[51][15].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane15_strm0_cntl          ( DownstreamStackBusLane[51][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane15_strm0_data          ( DownstreamStackBusLane[51][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane15_strm0_data_valid    ( DownstreamStackBusLane[51][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane15_strm1_ready         ( DownstreamStackBusLane[51][15].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane15_strm1_cntl          ( DownstreamStackBusLane[51][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane15_strm1_data          ( DownstreamStackBusLane[51][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane15_strm1_data_valid    ( DownstreamStackBusLane[51][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane16_strm0_ready         ( DownstreamStackBusLane[51][16].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane16_strm0_cntl          ( DownstreamStackBusLane[51][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane16_strm0_data          ( DownstreamStackBusLane[51][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane16_strm0_data_valid    ( DownstreamStackBusLane[51][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane16_strm1_ready         ( DownstreamStackBusLane[51][16].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane16_strm1_cntl          ( DownstreamStackBusLane[51][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane16_strm1_data          ( DownstreamStackBusLane[51][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane16_strm1_data_valid    ( DownstreamStackBusLane[51][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane17_strm0_ready         ( DownstreamStackBusLane[51][17].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane17_strm0_cntl          ( DownstreamStackBusLane[51][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane17_strm0_data          ( DownstreamStackBusLane[51][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane17_strm0_data_valid    ( DownstreamStackBusLane[51][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane17_strm1_ready         ( DownstreamStackBusLane[51][17].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane17_strm1_cntl          ( DownstreamStackBusLane[51][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane17_strm1_data          ( DownstreamStackBusLane[51][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane17_strm1_data_valid    ( DownstreamStackBusLane[51][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane18_strm0_ready         ( DownstreamStackBusLane[51][18].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane18_strm0_cntl          ( DownstreamStackBusLane[51][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane18_strm0_data          ( DownstreamStackBusLane[51][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane18_strm0_data_valid    ( DownstreamStackBusLane[51][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane18_strm1_ready         ( DownstreamStackBusLane[51][18].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane18_strm1_cntl          ( DownstreamStackBusLane[51][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane18_strm1_data          ( DownstreamStackBusLane[51][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane18_strm1_data_valid    ( DownstreamStackBusLane[51][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane19_strm0_ready         ( DownstreamStackBusLane[51][19].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane19_strm0_cntl          ( DownstreamStackBusLane[51][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane19_strm0_data          ( DownstreamStackBusLane[51][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane19_strm0_data_valid    ( DownstreamStackBusLane[51][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane19_strm1_ready         ( DownstreamStackBusLane[51][19].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane19_strm1_cntl          ( DownstreamStackBusLane[51][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane19_strm1_data          ( DownstreamStackBusLane[51][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane19_strm1_data_valid    ( DownstreamStackBusLane[51][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane20_strm0_ready         ( DownstreamStackBusLane[51][20].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane20_strm0_cntl          ( DownstreamStackBusLane[51][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane20_strm0_data          ( DownstreamStackBusLane[51][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane20_strm0_data_valid    ( DownstreamStackBusLane[51][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane20_strm1_ready         ( DownstreamStackBusLane[51][20].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane20_strm1_cntl          ( DownstreamStackBusLane[51][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane20_strm1_data          ( DownstreamStackBusLane[51][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane20_strm1_data_valid    ( DownstreamStackBusLane[51][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane21_strm0_ready         ( DownstreamStackBusLane[51][21].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane21_strm0_cntl          ( DownstreamStackBusLane[51][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane21_strm0_data          ( DownstreamStackBusLane[51][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane21_strm0_data_valid    ( DownstreamStackBusLane[51][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane21_strm1_ready         ( DownstreamStackBusLane[51][21].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane21_strm1_cntl          ( DownstreamStackBusLane[51][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane21_strm1_data          ( DownstreamStackBusLane[51][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane21_strm1_data_valid    ( DownstreamStackBusLane[51][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane22_strm0_ready         ( DownstreamStackBusLane[51][22].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane22_strm0_cntl          ( DownstreamStackBusLane[51][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane22_strm0_data          ( DownstreamStackBusLane[51][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane22_strm0_data_valid    ( DownstreamStackBusLane[51][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane22_strm1_ready         ( DownstreamStackBusLane[51][22].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane22_strm1_cntl          ( DownstreamStackBusLane[51][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane22_strm1_data          ( DownstreamStackBusLane[51][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane22_strm1_data_valid    ( DownstreamStackBusLane[51][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane23_strm0_ready         ( DownstreamStackBusLane[51][23].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane23_strm0_cntl          ( DownstreamStackBusLane[51][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane23_strm0_data          ( DownstreamStackBusLane[51][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane23_strm0_data_valid    ( DownstreamStackBusLane[51][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane23_strm1_ready         ( DownstreamStackBusLane[51][23].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane23_strm1_cntl          ( DownstreamStackBusLane[51][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane23_strm1_data          ( DownstreamStackBusLane[51][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane23_strm1_data_valid    ( DownstreamStackBusLane[51][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane24_strm0_ready         ( DownstreamStackBusLane[51][24].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane24_strm0_cntl          ( DownstreamStackBusLane[51][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane24_strm0_data          ( DownstreamStackBusLane[51][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane24_strm0_data_valid    ( DownstreamStackBusLane[51][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane24_strm1_ready         ( DownstreamStackBusLane[51][24].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane24_strm1_cntl          ( DownstreamStackBusLane[51][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane24_strm1_data          ( DownstreamStackBusLane[51][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane24_strm1_data_valid    ( DownstreamStackBusLane[51][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane25_strm0_ready         ( DownstreamStackBusLane[51][25].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane25_strm0_cntl          ( DownstreamStackBusLane[51][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane25_strm0_data          ( DownstreamStackBusLane[51][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane25_strm0_data_valid    ( DownstreamStackBusLane[51][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane25_strm1_ready         ( DownstreamStackBusLane[51][25].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane25_strm1_cntl          ( DownstreamStackBusLane[51][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane25_strm1_data          ( DownstreamStackBusLane[51][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane25_strm1_data_valid    ( DownstreamStackBusLane[51][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane26_strm0_ready         ( DownstreamStackBusLane[51][26].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane26_strm0_cntl          ( DownstreamStackBusLane[51][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane26_strm0_data          ( DownstreamStackBusLane[51][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane26_strm0_data_valid    ( DownstreamStackBusLane[51][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane26_strm1_ready         ( DownstreamStackBusLane[51][26].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane26_strm1_cntl          ( DownstreamStackBusLane[51][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane26_strm1_data          ( DownstreamStackBusLane[51][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane26_strm1_data_valid    ( DownstreamStackBusLane[51][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane27_strm0_ready         ( DownstreamStackBusLane[51][27].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane27_strm0_cntl          ( DownstreamStackBusLane[51][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane27_strm0_data          ( DownstreamStackBusLane[51][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane27_strm0_data_valid    ( DownstreamStackBusLane[51][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane27_strm1_ready         ( DownstreamStackBusLane[51][27].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane27_strm1_cntl          ( DownstreamStackBusLane[51][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane27_strm1_data          ( DownstreamStackBusLane[51][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane27_strm1_data_valid    ( DownstreamStackBusLane[51][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane28_strm0_ready         ( DownstreamStackBusLane[51][28].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane28_strm0_cntl          ( DownstreamStackBusLane[51][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane28_strm0_data          ( DownstreamStackBusLane[51][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane28_strm0_data_valid    ( DownstreamStackBusLane[51][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane28_strm1_ready         ( DownstreamStackBusLane[51][28].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane28_strm1_cntl          ( DownstreamStackBusLane[51][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane28_strm1_data          ( DownstreamStackBusLane[51][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane28_strm1_data_valid    ( DownstreamStackBusLane[51][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane29_strm0_ready         ( DownstreamStackBusLane[51][29].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane29_strm0_cntl          ( DownstreamStackBusLane[51][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane29_strm0_data          ( DownstreamStackBusLane[51][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane29_strm0_data_valid    ( DownstreamStackBusLane[51][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane29_strm1_ready         ( DownstreamStackBusLane[51][29].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane29_strm1_cntl          ( DownstreamStackBusLane[51][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane29_strm1_data          ( DownstreamStackBusLane[51][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane29_strm1_data_valid    ( DownstreamStackBusLane[51][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane30_strm0_ready         ( DownstreamStackBusLane[51][30].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane30_strm0_cntl          ( DownstreamStackBusLane[51][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane30_strm0_data          ( DownstreamStackBusLane[51][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane30_strm0_data_valid    ( DownstreamStackBusLane[51][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane30_strm1_ready         ( DownstreamStackBusLane[51][30].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane30_strm1_cntl          ( DownstreamStackBusLane[51][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane30_strm1_data          ( DownstreamStackBusLane[51][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane30_strm1_data_valid    ( DownstreamStackBusLane[51][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 51, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane31_strm0_ready         ( DownstreamStackBusLane[51][31].pe__std__lane_strm0_ready              ),      
        .std__pe51__lane31_strm0_cntl          ( DownstreamStackBusLane[51][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe51__lane31_strm0_data          ( DownstreamStackBusLane[51][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe51__lane31_strm0_data_valid    ( DownstreamStackBusLane[51][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__std__lane31_strm1_ready         ( DownstreamStackBusLane[51][31].pe__std__lane_strm1_ready              ),      
        .std__pe51__lane31_strm1_cntl          ( DownstreamStackBusLane[51][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe51__lane31_strm1_data          ( DownstreamStackBusLane[51][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe51__lane31_strm1_data_valid    ( DownstreamStackBusLane[51][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane0_strm0_ready         ( DownstreamStackBusLane[52][0].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane0_strm0_cntl          ( DownstreamStackBusLane[52][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane0_strm0_data          ( DownstreamStackBusLane[52][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane0_strm0_data_valid    ( DownstreamStackBusLane[52][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane0_strm1_ready         ( DownstreamStackBusLane[52][0].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane0_strm1_cntl          ( DownstreamStackBusLane[52][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane0_strm1_data          ( DownstreamStackBusLane[52][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane0_strm1_data_valid    ( DownstreamStackBusLane[52][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane1_strm0_ready         ( DownstreamStackBusLane[52][1].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane1_strm0_cntl          ( DownstreamStackBusLane[52][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane1_strm0_data          ( DownstreamStackBusLane[52][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane1_strm0_data_valid    ( DownstreamStackBusLane[52][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane1_strm1_ready         ( DownstreamStackBusLane[52][1].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane1_strm1_cntl          ( DownstreamStackBusLane[52][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane1_strm1_data          ( DownstreamStackBusLane[52][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane1_strm1_data_valid    ( DownstreamStackBusLane[52][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane2_strm0_ready         ( DownstreamStackBusLane[52][2].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane2_strm0_cntl          ( DownstreamStackBusLane[52][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane2_strm0_data          ( DownstreamStackBusLane[52][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane2_strm0_data_valid    ( DownstreamStackBusLane[52][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane2_strm1_ready         ( DownstreamStackBusLane[52][2].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane2_strm1_cntl          ( DownstreamStackBusLane[52][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane2_strm1_data          ( DownstreamStackBusLane[52][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane2_strm1_data_valid    ( DownstreamStackBusLane[52][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane3_strm0_ready         ( DownstreamStackBusLane[52][3].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane3_strm0_cntl          ( DownstreamStackBusLane[52][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane3_strm0_data          ( DownstreamStackBusLane[52][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane3_strm0_data_valid    ( DownstreamStackBusLane[52][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane3_strm1_ready         ( DownstreamStackBusLane[52][3].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane3_strm1_cntl          ( DownstreamStackBusLane[52][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane3_strm1_data          ( DownstreamStackBusLane[52][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane3_strm1_data_valid    ( DownstreamStackBusLane[52][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane4_strm0_ready         ( DownstreamStackBusLane[52][4].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane4_strm0_cntl          ( DownstreamStackBusLane[52][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane4_strm0_data          ( DownstreamStackBusLane[52][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane4_strm0_data_valid    ( DownstreamStackBusLane[52][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane4_strm1_ready         ( DownstreamStackBusLane[52][4].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane4_strm1_cntl          ( DownstreamStackBusLane[52][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane4_strm1_data          ( DownstreamStackBusLane[52][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane4_strm1_data_valid    ( DownstreamStackBusLane[52][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane5_strm0_ready         ( DownstreamStackBusLane[52][5].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane5_strm0_cntl          ( DownstreamStackBusLane[52][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane5_strm0_data          ( DownstreamStackBusLane[52][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane5_strm0_data_valid    ( DownstreamStackBusLane[52][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane5_strm1_ready         ( DownstreamStackBusLane[52][5].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane5_strm1_cntl          ( DownstreamStackBusLane[52][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane5_strm1_data          ( DownstreamStackBusLane[52][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane5_strm1_data_valid    ( DownstreamStackBusLane[52][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane6_strm0_ready         ( DownstreamStackBusLane[52][6].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane6_strm0_cntl          ( DownstreamStackBusLane[52][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane6_strm0_data          ( DownstreamStackBusLane[52][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane6_strm0_data_valid    ( DownstreamStackBusLane[52][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane6_strm1_ready         ( DownstreamStackBusLane[52][6].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane6_strm1_cntl          ( DownstreamStackBusLane[52][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane6_strm1_data          ( DownstreamStackBusLane[52][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane6_strm1_data_valid    ( DownstreamStackBusLane[52][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane7_strm0_ready         ( DownstreamStackBusLane[52][7].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane7_strm0_cntl          ( DownstreamStackBusLane[52][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane7_strm0_data          ( DownstreamStackBusLane[52][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane7_strm0_data_valid    ( DownstreamStackBusLane[52][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane7_strm1_ready         ( DownstreamStackBusLane[52][7].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane7_strm1_cntl          ( DownstreamStackBusLane[52][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane7_strm1_data          ( DownstreamStackBusLane[52][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane7_strm1_data_valid    ( DownstreamStackBusLane[52][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane8_strm0_ready         ( DownstreamStackBusLane[52][8].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane8_strm0_cntl          ( DownstreamStackBusLane[52][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane8_strm0_data          ( DownstreamStackBusLane[52][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane8_strm0_data_valid    ( DownstreamStackBusLane[52][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane8_strm1_ready         ( DownstreamStackBusLane[52][8].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane8_strm1_cntl          ( DownstreamStackBusLane[52][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane8_strm1_data          ( DownstreamStackBusLane[52][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane8_strm1_data_valid    ( DownstreamStackBusLane[52][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane9_strm0_ready         ( DownstreamStackBusLane[52][9].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane9_strm0_cntl          ( DownstreamStackBusLane[52][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane9_strm0_data          ( DownstreamStackBusLane[52][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane9_strm0_data_valid    ( DownstreamStackBusLane[52][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane9_strm1_ready         ( DownstreamStackBusLane[52][9].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane9_strm1_cntl          ( DownstreamStackBusLane[52][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane9_strm1_data          ( DownstreamStackBusLane[52][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane9_strm1_data_valid    ( DownstreamStackBusLane[52][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane10_strm0_ready         ( DownstreamStackBusLane[52][10].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane10_strm0_cntl          ( DownstreamStackBusLane[52][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane10_strm0_data          ( DownstreamStackBusLane[52][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane10_strm0_data_valid    ( DownstreamStackBusLane[52][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane10_strm1_ready         ( DownstreamStackBusLane[52][10].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane10_strm1_cntl          ( DownstreamStackBusLane[52][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane10_strm1_data          ( DownstreamStackBusLane[52][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane10_strm1_data_valid    ( DownstreamStackBusLane[52][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane11_strm0_ready         ( DownstreamStackBusLane[52][11].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane11_strm0_cntl          ( DownstreamStackBusLane[52][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane11_strm0_data          ( DownstreamStackBusLane[52][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane11_strm0_data_valid    ( DownstreamStackBusLane[52][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane11_strm1_ready         ( DownstreamStackBusLane[52][11].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane11_strm1_cntl          ( DownstreamStackBusLane[52][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane11_strm1_data          ( DownstreamStackBusLane[52][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane11_strm1_data_valid    ( DownstreamStackBusLane[52][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane12_strm0_ready         ( DownstreamStackBusLane[52][12].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane12_strm0_cntl          ( DownstreamStackBusLane[52][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane12_strm0_data          ( DownstreamStackBusLane[52][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane12_strm0_data_valid    ( DownstreamStackBusLane[52][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane12_strm1_ready         ( DownstreamStackBusLane[52][12].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane12_strm1_cntl          ( DownstreamStackBusLane[52][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane12_strm1_data          ( DownstreamStackBusLane[52][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane12_strm1_data_valid    ( DownstreamStackBusLane[52][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane13_strm0_ready         ( DownstreamStackBusLane[52][13].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane13_strm0_cntl          ( DownstreamStackBusLane[52][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane13_strm0_data          ( DownstreamStackBusLane[52][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane13_strm0_data_valid    ( DownstreamStackBusLane[52][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane13_strm1_ready         ( DownstreamStackBusLane[52][13].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane13_strm1_cntl          ( DownstreamStackBusLane[52][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane13_strm1_data          ( DownstreamStackBusLane[52][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane13_strm1_data_valid    ( DownstreamStackBusLane[52][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane14_strm0_ready         ( DownstreamStackBusLane[52][14].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane14_strm0_cntl          ( DownstreamStackBusLane[52][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane14_strm0_data          ( DownstreamStackBusLane[52][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane14_strm0_data_valid    ( DownstreamStackBusLane[52][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane14_strm1_ready         ( DownstreamStackBusLane[52][14].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane14_strm1_cntl          ( DownstreamStackBusLane[52][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane14_strm1_data          ( DownstreamStackBusLane[52][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane14_strm1_data_valid    ( DownstreamStackBusLane[52][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane15_strm0_ready         ( DownstreamStackBusLane[52][15].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane15_strm0_cntl          ( DownstreamStackBusLane[52][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane15_strm0_data          ( DownstreamStackBusLane[52][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane15_strm0_data_valid    ( DownstreamStackBusLane[52][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane15_strm1_ready         ( DownstreamStackBusLane[52][15].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane15_strm1_cntl          ( DownstreamStackBusLane[52][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane15_strm1_data          ( DownstreamStackBusLane[52][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane15_strm1_data_valid    ( DownstreamStackBusLane[52][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane16_strm0_ready         ( DownstreamStackBusLane[52][16].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane16_strm0_cntl          ( DownstreamStackBusLane[52][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane16_strm0_data          ( DownstreamStackBusLane[52][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane16_strm0_data_valid    ( DownstreamStackBusLane[52][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane16_strm1_ready         ( DownstreamStackBusLane[52][16].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane16_strm1_cntl          ( DownstreamStackBusLane[52][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane16_strm1_data          ( DownstreamStackBusLane[52][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane16_strm1_data_valid    ( DownstreamStackBusLane[52][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane17_strm0_ready         ( DownstreamStackBusLane[52][17].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane17_strm0_cntl          ( DownstreamStackBusLane[52][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane17_strm0_data          ( DownstreamStackBusLane[52][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane17_strm0_data_valid    ( DownstreamStackBusLane[52][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane17_strm1_ready         ( DownstreamStackBusLane[52][17].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane17_strm1_cntl          ( DownstreamStackBusLane[52][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane17_strm1_data          ( DownstreamStackBusLane[52][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane17_strm1_data_valid    ( DownstreamStackBusLane[52][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane18_strm0_ready         ( DownstreamStackBusLane[52][18].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane18_strm0_cntl          ( DownstreamStackBusLane[52][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane18_strm0_data          ( DownstreamStackBusLane[52][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane18_strm0_data_valid    ( DownstreamStackBusLane[52][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane18_strm1_ready         ( DownstreamStackBusLane[52][18].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane18_strm1_cntl          ( DownstreamStackBusLane[52][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane18_strm1_data          ( DownstreamStackBusLane[52][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane18_strm1_data_valid    ( DownstreamStackBusLane[52][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane19_strm0_ready         ( DownstreamStackBusLane[52][19].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane19_strm0_cntl          ( DownstreamStackBusLane[52][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane19_strm0_data          ( DownstreamStackBusLane[52][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane19_strm0_data_valid    ( DownstreamStackBusLane[52][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane19_strm1_ready         ( DownstreamStackBusLane[52][19].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane19_strm1_cntl          ( DownstreamStackBusLane[52][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane19_strm1_data          ( DownstreamStackBusLane[52][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane19_strm1_data_valid    ( DownstreamStackBusLane[52][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane20_strm0_ready         ( DownstreamStackBusLane[52][20].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane20_strm0_cntl          ( DownstreamStackBusLane[52][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane20_strm0_data          ( DownstreamStackBusLane[52][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane20_strm0_data_valid    ( DownstreamStackBusLane[52][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane20_strm1_ready         ( DownstreamStackBusLane[52][20].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane20_strm1_cntl          ( DownstreamStackBusLane[52][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane20_strm1_data          ( DownstreamStackBusLane[52][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane20_strm1_data_valid    ( DownstreamStackBusLane[52][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane21_strm0_ready         ( DownstreamStackBusLane[52][21].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane21_strm0_cntl          ( DownstreamStackBusLane[52][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane21_strm0_data          ( DownstreamStackBusLane[52][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane21_strm0_data_valid    ( DownstreamStackBusLane[52][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane21_strm1_ready         ( DownstreamStackBusLane[52][21].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane21_strm1_cntl          ( DownstreamStackBusLane[52][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane21_strm1_data          ( DownstreamStackBusLane[52][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane21_strm1_data_valid    ( DownstreamStackBusLane[52][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane22_strm0_ready         ( DownstreamStackBusLane[52][22].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane22_strm0_cntl          ( DownstreamStackBusLane[52][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane22_strm0_data          ( DownstreamStackBusLane[52][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane22_strm0_data_valid    ( DownstreamStackBusLane[52][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane22_strm1_ready         ( DownstreamStackBusLane[52][22].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane22_strm1_cntl          ( DownstreamStackBusLane[52][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane22_strm1_data          ( DownstreamStackBusLane[52][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane22_strm1_data_valid    ( DownstreamStackBusLane[52][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane23_strm0_ready         ( DownstreamStackBusLane[52][23].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane23_strm0_cntl          ( DownstreamStackBusLane[52][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane23_strm0_data          ( DownstreamStackBusLane[52][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane23_strm0_data_valid    ( DownstreamStackBusLane[52][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane23_strm1_ready         ( DownstreamStackBusLane[52][23].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane23_strm1_cntl          ( DownstreamStackBusLane[52][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane23_strm1_data          ( DownstreamStackBusLane[52][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane23_strm1_data_valid    ( DownstreamStackBusLane[52][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane24_strm0_ready         ( DownstreamStackBusLane[52][24].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane24_strm0_cntl          ( DownstreamStackBusLane[52][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane24_strm0_data          ( DownstreamStackBusLane[52][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane24_strm0_data_valid    ( DownstreamStackBusLane[52][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane24_strm1_ready         ( DownstreamStackBusLane[52][24].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane24_strm1_cntl          ( DownstreamStackBusLane[52][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane24_strm1_data          ( DownstreamStackBusLane[52][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane24_strm1_data_valid    ( DownstreamStackBusLane[52][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane25_strm0_ready         ( DownstreamStackBusLane[52][25].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane25_strm0_cntl          ( DownstreamStackBusLane[52][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane25_strm0_data          ( DownstreamStackBusLane[52][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane25_strm0_data_valid    ( DownstreamStackBusLane[52][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane25_strm1_ready         ( DownstreamStackBusLane[52][25].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane25_strm1_cntl          ( DownstreamStackBusLane[52][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane25_strm1_data          ( DownstreamStackBusLane[52][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane25_strm1_data_valid    ( DownstreamStackBusLane[52][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane26_strm0_ready         ( DownstreamStackBusLane[52][26].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane26_strm0_cntl          ( DownstreamStackBusLane[52][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane26_strm0_data          ( DownstreamStackBusLane[52][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane26_strm0_data_valid    ( DownstreamStackBusLane[52][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane26_strm1_ready         ( DownstreamStackBusLane[52][26].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane26_strm1_cntl          ( DownstreamStackBusLane[52][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane26_strm1_data          ( DownstreamStackBusLane[52][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane26_strm1_data_valid    ( DownstreamStackBusLane[52][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane27_strm0_ready         ( DownstreamStackBusLane[52][27].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane27_strm0_cntl          ( DownstreamStackBusLane[52][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane27_strm0_data          ( DownstreamStackBusLane[52][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane27_strm0_data_valid    ( DownstreamStackBusLane[52][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane27_strm1_ready         ( DownstreamStackBusLane[52][27].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane27_strm1_cntl          ( DownstreamStackBusLane[52][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane27_strm1_data          ( DownstreamStackBusLane[52][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane27_strm1_data_valid    ( DownstreamStackBusLane[52][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane28_strm0_ready         ( DownstreamStackBusLane[52][28].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane28_strm0_cntl          ( DownstreamStackBusLane[52][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane28_strm0_data          ( DownstreamStackBusLane[52][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane28_strm0_data_valid    ( DownstreamStackBusLane[52][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane28_strm1_ready         ( DownstreamStackBusLane[52][28].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane28_strm1_cntl          ( DownstreamStackBusLane[52][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane28_strm1_data          ( DownstreamStackBusLane[52][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane28_strm1_data_valid    ( DownstreamStackBusLane[52][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane29_strm0_ready         ( DownstreamStackBusLane[52][29].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane29_strm0_cntl          ( DownstreamStackBusLane[52][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane29_strm0_data          ( DownstreamStackBusLane[52][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane29_strm0_data_valid    ( DownstreamStackBusLane[52][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane29_strm1_ready         ( DownstreamStackBusLane[52][29].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane29_strm1_cntl          ( DownstreamStackBusLane[52][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane29_strm1_data          ( DownstreamStackBusLane[52][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane29_strm1_data_valid    ( DownstreamStackBusLane[52][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane30_strm0_ready         ( DownstreamStackBusLane[52][30].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane30_strm0_cntl          ( DownstreamStackBusLane[52][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane30_strm0_data          ( DownstreamStackBusLane[52][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane30_strm0_data_valid    ( DownstreamStackBusLane[52][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane30_strm1_ready         ( DownstreamStackBusLane[52][30].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane30_strm1_cntl          ( DownstreamStackBusLane[52][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane30_strm1_data          ( DownstreamStackBusLane[52][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane30_strm1_data_valid    ( DownstreamStackBusLane[52][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 52, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane31_strm0_ready         ( DownstreamStackBusLane[52][31].pe__std__lane_strm0_ready              ),      
        .std__pe52__lane31_strm0_cntl          ( DownstreamStackBusLane[52][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe52__lane31_strm0_data          ( DownstreamStackBusLane[52][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe52__lane31_strm0_data_valid    ( DownstreamStackBusLane[52][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__std__lane31_strm1_ready         ( DownstreamStackBusLane[52][31].pe__std__lane_strm1_ready              ),      
        .std__pe52__lane31_strm1_cntl          ( DownstreamStackBusLane[52][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe52__lane31_strm1_data          ( DownstreamStackBusLane[52][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe52__lane31_strm1_data_valid    ( DownstreamStackBusLane[52][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane0_strm0_ready         ( DownstreamStackBusLane[53][0].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane0_strm0_cntl          ( DownstreamStackBusLane[53][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane0_strm0_data          ( DownstreamStackBusLane[53][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane0_strm0_data_valid    ( DownstreamStackBusLane[53][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane0_strm1_ready         ( DownstreamStackBusLane[53][0].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane0_strm1_cntl          ( DownstreamStackBusLane[53][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane0_strm1_data          ( DownstreamStackBusLane[53][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane0_strm1_data_valid    ( DownstreamStackBusLane[53][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane1_strm0_ready         ( DownstreamStackBusLane[53][1].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane1_strm0_cntl          ( DownstreamStackBusLane[53][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane1_strm0_data          ( DownstreamStackBusLane[53][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane1_strm0_data_valid    ( DownstreamStackBusLane[53][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane1_strm1_ready         ( DownstreamStackBusLane[53][1].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane1_strm1_cntl          ( DownstreamStackBusLane[53][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane1_strm1_data          ( DownstreamStackBusLane[53][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane1_strm1_data_valid    ( DownstreamStackBusLane[53][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane2_strm0_ready         ( DownstreamStackBusLane[53][2].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane2_strm0_cntl          ( DownstreamStackBusLane[53][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane2_strm0_data          ( DownstreamStackBusLane[53][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane2_strm0_data_valid    ( DownstreamStackBusLane[53][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane2_strm1_ready         ( DownstreamStackBusLane[53][2].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane2_strm1_cntl          ( DownstreamStackBusLane[53][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane2_strm1_data          ( DownstreamStackBusLane[53][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane2_strm1_data_valid    ( DownstreamStackBusLane[53][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane3_strm0_ready         ( DownstreamStackBusLane[53][3].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane3_strm0_cntl          ( DownstreamStackBusLane[53][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane3_strm0_data          ( DownstreamStackBusLane[53][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane3_strm0_data_valid    ( DownstreamStackBusLane[53][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane3_strm1_ready         ( DownstreamStackBusLane[53][3].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane3_strm1_cntl          ( DownstreamStackBusLane[53][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane3_strm1_data          ( DownstreamStackBusLane[53][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane3_strm1_data_valid    ( DownstreamStackBusLane[53][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane4_strm0_ready         ( DownstreamStackBusLane[53][4].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane4_strm0_cntl          ( DownstreamStackBusLane[53][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane4_strm0_data          ( DownstreamStackBusLane[53][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane4_strm0_data_valid    ( DownstreamStackBusLane[53][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane4_strm1_ready         ( DownstreamStackBusLane[53][4].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane4_strm1_cntl          ( DownstreamStackBusLane[53][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane4_strm1_data          ( DownstreamStackBusLane[53][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane4_strm1_data_valid    ( DownstreamStackBusLane[53][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane5_strm0_ready         ( DownstreamStackBusLane[53][5].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane5_strm0_cntl          ( DownstreamStackBusLane[53][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane5_strm0_data          ( DownstreamStackBusLane[53][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane5_strm0_data_valid    ( DownstreamStackBusLane[53][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane5_strm1_ready         ( DownstreamStackBusLane[53][5].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane5_strm1_cntl          ( DownstreamStackBusLane[53][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane5_strm1_data          ( DownstreamStackBusLane[53][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane5_strm1_data_valid    ( DownstreamStackBusLane[53][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane6_strm0_ready         ( DownstreamStackBusLane[53][6].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane6_strm0_cntl          ( DownstreamStackBusLane[53][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane6_strm0_data          ( DownstreamStackBusLane[53][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane6_strm0_data_valid    ( DownstreamStackBusLane[53][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane6_strm1_ready         ( DownstreamStackBusLane[53][6].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane6_strm1_cntl          ( DownstreamStackBusLane[53][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane6_strm1_data          ( DownstreamStackBusLane[53][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane6_strm1_data_valid    ( DownstreamStackBusLane[53][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane7_strm0_ready         ( DownstreamStackBusLane[53][7].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane7_strm0_cntl          ( DownstreamStackBusLane[53][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane7_strm0_data          ( DownstreamStackBusLane[53][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane7_strm0_data_valid    ( DownstreamStackBusLane[53][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane7_strm1_ready         ( DownstreamStackBusLane[53][7].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane7_strm1_cntl          ( DownstreamStackBusLane[53][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane7_strm1_data          ( DownstreamStackBusLane[53][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane7_strm1_data_valid    ( DownstreamStackBusLane[53][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane8_strm0_ready         ( DownstreamStackBusLane[53][8].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane8_strm0_cntl          ( DownstreamStackBusLane[53][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane8_strm0_data          ( DownstreamStackBusLane[53][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane8_strm0_data_valid    ( DownstreamStackBusLane[53][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane8_strm1_ready         ( DownstreamStackBusLane[53][8].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane8_strm1_cntl          ( DownstreamStackBusLane[53][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane8_strm1_data          ( DownstreamStackBusLane[53][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane8_strm1_data_valid    ( DownstreamStackBusLane[53][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane9_strm0_ready         ( DownstreamStackBusLane[53][9].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane9_strm0_cntl          ( DownstreamStackBusLane[53][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane9_strm0_data          ( DownstreamStackBusLane[53][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane9_strm0_data_valid    ( DownstreamStackBusLane[53][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane9_strm1_ready         ( DownstreamStackBusLane[53][9].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane9_strm1_cntl          ( DownstreamStackBusLane[53][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane9_strm1_data          ( DownstreamStackBusLane[53][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane9_strm1_data_valid    ( DownstreamStackBusLane[53][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane10_strm0_ready         ( DownstreamStackBusLane[53][10].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane10_strm0_cntl          ( DownstreamStackBusLane[53][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane10_strm0_data          ( DownstreamStackBusLane[53][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane10_strm0_data_valid    ( DownstreamStackBusLane[53][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane10_strm1_ready         ( DownstreamStackBusLane[53][10].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane10_strm1_cntl          ( DownstreamStackBusLane[53][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane10_strm1_data          ( DownstreamStackBusLane[53][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane10_strm1_data_valid    ( DownstreamStackBusLane[53][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane11_strm0_ready         ( DownstreamStackBusLane[53][11].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane11_strm0_cntl          ( DownstreamStackBusLane[53][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane11_strm0_data          ( DownstreamStackBusLane[53][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane11_strm0_data_valid    ( DownstreamStackBusLane[53][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane11_strm1_ready         ( DownstreamStackBusLane[53][11].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane11_strm1_cntl          ( DownstreamStackBusLane[53][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane11_strm1_data          ( DownstreamStackBusLane[53][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane11_strm1_data_valid    ( DownstreamStackBusLane[53][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane12_strm0_ready         ( DownstreamStackBusLane[53][12].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane12_strm0_cntl          ( DownstreamStackBusLane[53][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane12_strm0_data          ( DownstreamStackBusLane[53][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane12_strm0_data_valid    ( DownstreamStackBusLane[53][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane12_strm1_ready         ( DownstreamStackBusLane[53][12].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane12_strm1_cntl          ( DownstreamStackBusLane[53][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane12_strm1_data          ( DownstreamStackBusLane[53][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane12_strm1_data_valid    ( DownstreamStackBusLane[53][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane13_strm0_ready         ( DownstreamStackBusLane[53][13].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane13_strm0_cntl          ( DownstreamStackBusLane[53][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane13_strm0_data          ( DownstreamStackBusLane[53][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane13_strm0_data_valid    ( DownstreamStackBusLane[53][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane13_strm1_ready         ( DownstreamStackBusLane[53][13].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane13_strm1_cntl          ( DownstreamStackBusLane[53][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane13_strm1_data          ( DownstreamStackBusLane[53][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane13_strm1_data_valid    ( DownstreamStackBusLane[53][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane14_strm0_ready         ( DownstreamStackBusLane[53][14].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane14_strm0_cntl          ( DownstreamStackBusLane[53][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane14_strm0_data          ( DownstreamStackBusLane[53][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane14_strm0_data_valid    ( DownstreamStackBusLane[53][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane14_strm1_ready         ( DownstreamStackBusLane[53][14].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane14_strm1_cntl          ( DownstreamStackBusLane[53][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane14_strm1_data          ( DownstreamStackBusLane[53][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane14_strm1_data_valid    ( DownstreamStackBusLane[53][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane15_strm0_ready         ( DownstreamStackBusLane[53][15].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane15_strm0_cntl          ( DownstreamStackBusLane[53][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane15_strm0_data          ( DownstreamStackBusLane[53][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane15_strm0_data_valid    ( DownstreamStackBusLane[53][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane15_strm1_ready         ( DownstreamStackBusLane[53][15].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane15_strm1_cntl          ( DownstreamStackBusLane[53][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane15_strm1_data          ( DownstreamStackBusLane[53][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane15_strm1_data_valid    ( DownstreamStackBusLane[53][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane16_strm0_ready         ( DownstreamStackBusLane[53][16].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane16_strm0_cntl          ( DownstreamStackBusLane[53][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane16_strm0_data          ( DownstreamStackBusLane[53][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane16_strm0_data_valid    ( DownstreamStackBusLane[53][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane16_strm1_ready         ( DownstreamStackBusLane[53][16].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane16_strm1_cntl          ( DownstreamStackBusLane[53][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane16_strm1_data          ( DownstreamStackBusLane[53][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane16_strm1_data_valid    ( DownstreamStackBusLane[53][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane17_strm0_ready         ( DownstreamStackBusLane[53][17].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane17_strm0_cntl          ( DownstreamStackBusLane[53][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane17_strm0_data          ( DownstreamStackBusLane[53][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane17_strm0_data_valid    ( DownstreamStackBusLane[53][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane17_strm1_ready         ( DownstreamStackBusLane[53][17].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane17_strm1_cntl          ( DownstreamStackBusLane[53][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane17_strm1_data          ( DownstreamStackBusLane[53][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane17_strm1_data_valid    ( DownstreamStackBusLane[53][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane18_strm0_ready         ( DownstreamStackBusLane[53][18].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane18_strm0_cntl          ( DownstreamStackBusLane[53][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane18_strm0_data          ( DownstreamStackBusLane[53][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane18_strm0_data_valid    ( DownstreamStackBusLane[53][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane18_strm1_ready         ( DownstreamStackBusLane[53][18].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane18_strm1_cntl          ( DownstreamStackBusLane[53][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane18_strm1_data          ( DownstreamStackBusLane[53][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane18_strm1_data_valid    ( DownstreamStackBusLane[53][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane19_strm0_ready         ( DownstreamStackBusLane[53][19].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane19_strm0_cntl          ( DownstreamStackBusLane[53][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane19_strm0_data          ( DownstreamStackBusLane[53][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane19_strm0_data_valid    ( DownstreamStackBusLane[53][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane19_strm1_ready         ( DownstreamStackBusLane[53][19].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane19_strm1_cntl          ( DownstreamStackBusLane[53][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane19_strm1_data          ( DownstreamStackBusLane[53][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane19_strm1_data_valid    ( DownstreamStackBusLane[53][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane20_strm0_ready         ( DownstreamStackBusLane[53][20].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane20_strm0_cntl          ( DownstreamStackBusLane[53][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane20_strm0_data          ( DownstreamStackBusLane[53][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane20_strm0_data_valid    ( DownstreamStackBusLane[53][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane20_strm1_ready         ( DownstreamStackBusLane[53][20].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane20_strm1_cntl          ( DownstreamStackBusLane[53][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane20_strm1_data          ( DownstreamStackBusLane[53][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane20_strm1_data_valid    ( DownstreamStackBusLane[53][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane21_strm0_ready         ( DownstreamStackBusLane[53][21].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane21_strm0_cntl          ( DownstreamStackBusLane[53][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane21_strm0_data          ( DownstreamStackBusLane[53][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane21_strm0_data_valid    ( DownstreamStackBusLane[53][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane21_strm1_ready         ( DownstreamStackBusLane[53][21].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane21_strm1_cntl          ( DownstreamStackBusLane[53][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane21_strm1_data          ( DownstreamStackBusLane[53][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane21_strm1_data_valid    ( DownstreamStackBusLane[53][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane22_strm0_ready         ( DownstreamStackBusLane[53][22].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane22_strm0_cntl          ( DownstreamStackBusLane[53][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane22_strm0_data          ( DownstreamStackBusLane[53][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane22_strm0_data_valid    ( DownstreamStackBusLane[53][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane22_strm1_ready         ( DownstreamStackBusLane[53][22].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane22_strm1_cntl          ( DownstreamStackBusLane[53][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane22_strm1_data          ( DownstreamStackBusLane[53][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane22_strm1_data_valid    ( DownstreamStackBusLane[53][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane23_strm0_ready         ( DownstreamStackBusLane[53][23].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane23_strm0_cntl          ( DownstreamStackBusLane[53][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane23_strm0_data          ( DownstreamStackBusLane[53][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane23_strm0_data_valid    ( DownstreamStackBusLane[53][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane23_strm1_ready         ( DownstreamStackBusLane[53][23].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane23_strm1_cntl          ( DownstreamStackBusLane[53][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane23_strm1_data          ( DownstreamStackBusLane[53][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane23_strm1_data_valid    ( DownstreamStackBusLane[53][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane24_strm0_ready         ( DownstreamStackBusLane[53][24].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane24_strm0_cntl          ( DownstreamStackBusLane[53][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane24_strm0_data          ( DownstreamStackBusLane[53][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane24_strm0_data_valid    ( DownstreamStackBusLane[53][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane24_strm1_ready         ( DownstreamStackBusLane[53][24].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane24_strm1_cntl          ( DownstreamStackBusLane[53][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane24_strm1_data          ( DownstreamStackBusLane[53][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane24_strm1_data_valid    ( DownstreamStackBusLane[53][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane25_strm0_ready         ( DownstreamStackBusLane[53][25].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane25_strm0_cntl          ( DownstreamStackBusLane[53][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane25_strm0_data          ( DownstreamStackBusLane[53][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane25_strm0_data_valid    ( DownstreamStackBusLane[53][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane25_strm1_ready         ( DownstreamStackBusLane[53][25].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane25_strm1_cntl          ( DownstreamStackBusLane[53][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane25_strm1_data          ( DownstreamStackBusLane[53][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane25_strm1_data_valid    ( DownstreamStackBusLane[53][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane26_strm0_ready         ( DownstreamStackBusLane[53][26].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane26_strm0_cntl          ( DownstreamStackBusLane[53][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane26_strm0_data          ( DownstreamStackBusLane[53][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane26_strm0_data_valid    ( DownstreamStackBusLane[53][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane26_strm1_ready         ( DownstreamStackBusLane[53][26].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane26_strm1_cntl          ( DownstreamStackBusLane[53][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane26_strm1_data          ( DownstreamStackBusLane[53][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane26_strm1_data_valid    ( DownstreamStackBusLane[53][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane27_strm0_ready         ( DownstreamStackBusLane[53][27].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane27_strm0_cntl          ( DownstreamStackBusLane[53][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane27_strm0_data          ( DownstreamStackBusLane[53][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane27_strm0_data_valid    ( DownstreamStackBusLane[53][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane27_strm1_ready         ( DownstreamStackBusLane[53][27].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane27_strm1_cntl          ( DownstreamStackBusLane[53][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane27_strm1_data          ( DownstreamStackBusLane[53][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane27_strm1_data_valid    ( DownstreamStackBusLane[53][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane28_strm0_ready         ( DownstreamStackBusLane[53][28].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane28_strm0_cntl          ( DownstreamStackBusLane[53][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane28_strm0_data          ( DownstreamStackBusLane[53][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane28_strm0_data_valid    ( DownstreamStackBusLane[53][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane28_strm1_ready         ( DownstreamStackBusLane[53][28].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane28_strm1_cntl          ( DownstreamStackBusLane[53][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane28_strm1_data          ( DownstreamStackBusLane[53][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane28_strm1_data_valid    ( DownstreamStackBusLane[53][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane29_strm0_ready         ( DownstreamStackBusLane[53][29].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane29_strm0_cntl          ( DownstreamStackBusLane[53][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane29_strm0_data          ( DownstreamStackBusLane[53][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane29_strm0_data_valid    ( DownstreamStackBusLane[53][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane29_strm1_ready         ( DownstreamStackBusLane[53][29].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane29_strm1_cntl          ( DownstreamStackBusLane[53][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane29_strm1_data          ( DownstreamStackBusLane[53][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane29_strm1_data_valid    ( DownstreamStackBusLane[53][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane30_strm0_ready         ( DownstreamStackBusLane[53][30].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane30_strm0_cntl          ( DownstreamStackBusLane[53][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane30_strm0_data          ( DownstreamStackBusLane[53][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane30_strm0_data_valid    ( DownstreamStackBusLane[53][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane30_strm1_ready         ( DownstreamStackBusLane[53][30].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane30_strm1_cntl          ( DownstreamStackBusLane[53][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane30_strm1_data          ( DownstreamStackBusLane[53][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane30_strm1_data_valid    ( DownstreamStackBusLane[53][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 53, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane31_strm0_ready         ( DownstreamStackBusLane[53][31].pe__std__lane_strm0_ready              ),      
        .std__pe53__lane31_strm0_cntl          ( DownstreamStackBusLane[53][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe53__lane31_strm0_data          ( DownstreamStackBusLane[53][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe53__lane31_strm0_data_valid    ( DownstreamStackBusLane[53][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__std__lane31_strm1_ready         ( DownstreamStackBusLane[53][31].pe__std__lane_strm1_ready              ),      
        .std__pe53__lane31_strm1_cntl          ( DownstreamStackBusLane[53][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe53__lane31_strm1_data          ( DownstreamStackBusLane[53][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe53__lane31_strm1_data_valid    ( DownstreamStackBusLane[53][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane0_strm0_ready         ( DownstreamStackBusLane[54][0].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane0_strm0_cntl          ( DownstreamStackBusLane[54][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane0_strm0_data          ( DownstreamStackBusLane[54][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane0_strm0_data_valid    ( DownstreamStackBusLane[54][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane0_strm1_ready         ( DownstreamStackBusLane[54][0].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane0_strm1_cntl          ( DownstreamStackBusLane[54][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane0_strm1_data          ( DownstreamStackBusLane[54][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane0_strm1_data_valid    ( DownstreamStackBusLane[54][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane1_strm0_ready         ( DownstreamStackBusLane[54][1].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane1_strm0_cntl          ( DownstreamStackBusLane[54][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane1_strm0_data          ( DownstreamStackBusLane[54][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane1_strm0_data_valid    ( DownstreamStackBusLane[54][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane1_strm1_ready         ( DownstreamStackBusLane[54][1].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane1_strm1_cntl          ( DownstreamStackBusLane[54][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane1_strm1_data          ( DownstreamStackBusLane[54][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane1_strm1_data_valid    ( DownstreamStackBusLane[54][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane2_strm0_ready         ( DownstreamStackBusLane[54][2].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane2_strm0_cntl          ( DownstreamStackBusLane[54][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane2_strm0_data          ( DownstreamStackBusLane[54][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane2_strm0_data_valid    ( DownstreamStackBusLane[54][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane2_strm1_ready         ( DownstreamStackBusLane[54][2].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane2_strm1_cntl          ( DownstreamStackBusLane[54][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane2_strm1_data          ( DownstreamStackBusLane[54][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane2_strm1_data_valid    ( DownstreamStackBusLane[54][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane3_strm0_ready         ( DownstreamStackBusLane[54][3].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane3_strm0_cntl          ( DownstreamStackBusLane[54][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane3_strm0_data          ( DownstreamStackBusLane[54][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane3_strm0_data_valid    ( DownstreamStackBusLane[54][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane3_strm1_ready         ( DownstreamStackBusLane[54][3].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane3_strm1_cntl          ( DownstreamStackBusLane[54][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane3_strm1_data          ( DownstreamStackBusLane[54][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane3_strm1_data_valid    ( DownstreamStackBusLane[54][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane4_strm0_ready         ( DownstreamStackBusLane[54][4].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane4_strm0_cntl          ( DownstreamStackBusLane[54][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane4_strm0_data          ( DownstreamStackBusLane[54][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane4_strm0_data_valid    ( DownstreamStackBusLane[54][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane4_strm1_ready         ( DownstreamStackBusLane[54][4].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane4_strm1_cntl          ( DownstreamStackBusLane[54][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane4_strm1_data          ( DownstreamStackBusLane[54][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane4_strm1_data_valid    ( DownstreamStackBusLane[54][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane5_strm0_ready         ( DownstreamStackBusLane[54][5].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane5_strm0_cntl          ( DownstreamStackBusLane[54][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane5_strm0_data          ( DownstreamStackBusLane[54][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane5_strm0_data_valid    ( DownstreamStackBusLane[54][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane5_strm1_ready         ( DownstreamStackBusLane[54][5].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane5_strm1_cntl          ( DownstreamStackBusLane[54][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane5_strm1_data          ( DownstreamStackBusLane[54][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane5_strm1_data_valid    ( DownstreamStackBusLane[54][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane6_strm0_ready         ( DownstreamStackBusLane[54][6].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane6_strm0_cntl          ( DownstreamStackBusLane[54][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane6_strm0_data          ( DownstreamStackBusLane[54][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane6_strm0_data_valid    ( DownstreamStackBusLane[54][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane6_strm1_ready         ( DownstreamStackBusLane[54][6].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane6_strm1_cntl          ( DownstreamStackBusLane[54][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane6_strm1_data          ( DownstreamStackBusLane[54][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane6_strm1_data_valid    ( DownstreamStackBusLane[54][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane7_strm0_ready         ( DownstreamStackBusLane[54][7].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane7_strm0_cntl          ( DownstreamStackBusLane[54][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane7_strm0_data          ( DownstreamStackBusLane[54][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane7_strm0_data_valid    ( DownstreamStackBusLane[54][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane7_strm1_ready         ( DownstreamStackBusLane[54][7].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane7_strm1_cntl          ( DownstreamStackBusLane[54][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane7_strm1_data          ( DownstreamStackBusLane[54][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane7_strm1_data_valid    ( DownstreamStackBusLane[54][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane8_strm0_ready         ( DownstreamStackBusLane[54][8].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane8_strm0_cntl          ( DownstreamStackBusLane[54][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane8_strm0_data          ( DownstreamStackBusLane[54][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane8_strm0_data_valid    ( DownstreamStackBusLane[54][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane8_strm1_ready         ( DownstreamStackBusLane[54][8].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane8_strm1_cntl          ( DownstreamStackBusLane[54][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane8_strm1_data          ( DownstreamStackBusLane[54][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane8_strm1_data_valid    ( DownstreamStackBusLane[54][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane9_strm0_ready         ( DownstreamStackBusLane[54][9].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane9_strm0_cntl          ( DownstreamStackBusLane[54][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane9_strm0_data          ( DownstreamStackBusLane[54][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane9_strm0_data_valid    ( DownstreamStackBusLane[54][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane9_strm1_ready         ( DownstreamStackBusLane[54][9].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane9_strm1_cntl          ( DownstreamStackBusLane[54][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane9_strm1_data          ( DownstreamStackBusLane[54][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane9_strm1_data_valid    ( DownstreamStackBusLane[54][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane10_strm0_ready         ( DownstreamStackBusLane[54][10].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane10_strm0_cntl          ( DownstreamStackBusLane[54][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane10_strm0_data          ( DownstreamStackBusLane[54][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane10_strm0_data_valid    ( DownstreamStackBusLane[54][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane10_strm1_ready         ( DownstreamStackBusLane[54][10].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane10_strm1_cntl          ( DownstreamStackBusLane[54][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane10_strm1_data          ( DownstreamStackBusLane[54][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane10_strm1_data_valid    ( DownstreamStackBusLane[54][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane11_strm0_ready         ( DownstreamStackBusLane[54][11].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane11_strm0_cntl          ( DownstreamStackBusLane[54][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane11_strm0_data          ( DownstreamStackBusLane[54][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane11_strm0_data_valid    ( DownstreamStackBusLane[54][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane11_strm1_ready         ( DownstreamStackBusLane[54][11].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane11_strm1_cntl          ( DownstreamStackBusLane[54][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane11_strm1_data          ( DownstreamStackBusLane[54][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane11_strm1_data_valid    ( DownstreamStackBusLane[54][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane12_strm0_ready         ( DownstreamStackBusLane[54][12].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane12_strm0_cntl          ( DownstreamStackBusLane[54][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane12_strm0_data          ( DownstreamStackBusLane[54][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane12_strm0_data_valid    ( DownstreamStackBusLane[54][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane12_strm1_ready         ( DownstreamStackBusLane[54][12].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane12_strm1_cntl          ( DownstreamStackBusLane[54][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane12_strm1_data          ( DownstreamStackBusLane[54][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane12_strm1_data_valid    ( DownstreamStackBusLane[54][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane13_strm0_ready         ( DownstreamStackBusLane[54][13].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane13_strm0_cntl          ( DownstreamStackBusLane[54][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane13_strm0_data          ( DownstreamStackBusLane[54][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane13_strm0_data_valid    ( DownstreamStackBusLane[54][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane13_strm1_ready         ( DownstreamStackBusLane[54][13].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane13_strm1_cntl          ( DownstreamStackBusLane[54][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane13_strm1_data          ( DownstreamStackBusLane[54][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane13_strm1_data_valid    ( DownstreamStackBusLane[54][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane14_strm0_ready         ( DownstreamStackBusLane[54][14].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane14_strm0_cntl          ( DownstreamStackBusLane[54][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane14_strm0_data          ( DownstreamStackBusLane[54][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane14_strm0_data_valid    ( DownstreamStackBusLane[54][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane14_strm1_ready         ( DownstreamStackBusLane[54][14].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane14_strm1_cntl          ( DownstreamStackBusLane[54][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane14_strm1_data          ( DownstreamStackBusLane[54][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane14_strm1_data_valid    ( DownstreamStackBusLane[54][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane15_strm0_ready         ( DownstreamStackBusLane[54][15].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane15_strm0_cntl          ( DownstreamStackBusLane[54][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane15_strm0_data          ( DownstreamStackBusLane[54][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane15_strm0_data_valid    ( DownstreamStackBusLane[54][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane15_strm1_ready         ( DownstreamStackBusLane[54][15].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane15_strm1_cntl          ( DownstreamStackBusLane[54][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane15_strm1_data          ( DownstreamStackBusLane[54][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane15_strm1_data_valid    ( DownstreamStackBusLane[54][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane16_strm0_ready         ( DownstreamStackBusLane[54][16].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane16_strm0_cntl          ( DownstreamStackBusLane[54][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane16_strm0_data          ( DownstreamStackBusLane[54][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane16_strm0_data_valid    ( DownstreamStackBusLane[54][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane16_strm1_ready         ( DownstreamStackBusLane[54][16].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane16_strm1_cntl          ( DownstreamStackBusLane[54][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane16_strm1_data          ( DownstreamStackBusLane[54][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane16_strm1_data_valid    ( DownstreamStackBusLane[54][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane17_strm0_ready         ( DownstreamStackBusLane[54][17].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane17_strm0_cntl          ( DownstreamStackBusLane[54][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane17_strm0_data          ( DownstreamStackBusLane[54][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane17_strm0_data_valid    ( DownstreamStackBusLane[54][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane17_strm1_ready         ( DownstreamStackBusLane[54][17].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane17_strm1_cntl          ( DownstreamStackBusLane[54][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane17_strm1_data          ( DownstreamStackBusLane[54][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane17_strm1_data_valid    ( DownstreamStackBusLane[54][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane18_strm0_ready         ( DownstreamStackBusLane[54][18].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane18_strm0_cntl          ( DownstreamStackBusLane[54][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane18_strm0_data          ( DownstreamStackBusLane[54][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane18_strm0_data_valid    ( DownstreamStackBusLane[54][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane18_strm1_ready         ( DownstreamStackBusLane[54][18].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane18_strm1_cntl          ( DownstreamStackBusLane[54][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane18_strm1_data          ( DownstreamStackBusLane[54][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane18_strm1_data_valid    ( DownstreamStackBusLane[54][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane19_strm0_ready         ( DownstreamStackBusLane[54][19].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane19_strm0_cntl          ( DownstreamStackBusLane[54][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane19_strm0_data          ( DownstreamStackBusLane[54][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane19_strm0_data_valid    ( DownstreamStackBusLane[54][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane19_strm1_ready         ( DownstreamStackBusLane[54][19].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane19_strm1_cntl          ( DownstreamStackBusLane[54][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane19_strm1_data          ( DownstreamStackBusLane[54][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane19_strm1_data_valid    ( DownstreamStackBusLane[54][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane20_strm0_ready         ( DownstreamStackBusLane[54][20].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane20_strm0_cntl          ( DownstreamStackBusLane[54][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane20_strm0_data          ( DownstreamStackBusLane[54][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane20_strm0_data_valid    ( DownstreamStackBusLane[54][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane20_strm1_ready         ( DownstreamStackBusLane[54][20].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane20_strm1_cntl          ( DownstreamStackBusLane[54][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane20_strm1_data          ( DownstreamStackBusLane[54][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane20_strm1_data_valid    ( DownstreamStackBusLane[54][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane21_strm0_ready         ( DownstreamStackBusLane[54][21].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane21_strm0_cntl          ( DownstreamStackBusLane[54][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane21_strm0_data          ( DownstreamStackBusLane[54][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane21_strm0_data_valid    ( DownstreamStackBusLane[54][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane21_strm1_ready         ( DownstreamStackBusLane[54][21].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane21_strm1_cntl          ( DownstreamStackBusLane[54][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane21_strm1_data          ( DownstreamStackBusLane[54][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane21_strm1_data_valid    ( DownstreamStackBusLane[54][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane22_strm0_ready         ( DownstreamStackBusLane[54][22].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane22_strm0_cntl          ( DownstreamStackBusLane[54][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane22_strm0_data          ( DownstreamStackBusLane[54][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane22_strm0_data_valid    ( DownstreamStackBusLane[54][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane22_strm1_ready         ( DownstreamStackBusLane[54][22].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane22_strm1_cntl          ( DownstreamStackBusLane[54][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane22_strm1_data          ( DownstreamStackBusLane[54][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane22_strm1_data_valid    ( DownstreamStackBusLane[54][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane23_strm0_ready         ( DownstreamStackBusLane[54][23].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane23_strm0_cntl          ( DownstreamStackBusLane[54][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane23_strm0_data          ( DownstreamStackBusLane[54][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane23_strm0_data_valid    ( DownstreamStackBusLane[54][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane23_strm1_ready         ( DownstreamStackBusLane[54][23].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane23_strm1_cntl          ( DownstreamStackBusLane[54][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane23_strm1_data          ( DownstreamStackBusLane[54][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane23_strm1_data_valid    ( DownstreamStackBusLane[54][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane24_strm0_ready         ( DownstreamStackBusLane[54][24].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane24_strm0_cntl          ( DownstreamStackBusLane[54][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane24_strm0_data          ( DownstreamStackBusLane[54][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane24_strm0_data_valid    ( DownstreamStackBusLane[54][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane24_strm1_ready         ( DownstreamStackBusLane[54][24].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane24_strm1_cntl          ( DownstreamStackBusLane[54][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane24_strm1_data          ( DownstreamStackBusLane[54][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane24_strm1_data_valid    ( DownstreamStackBusLane[54][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane25_strm0_ready         ( DownstreamStackBusLane[54][25].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane25_strm0_cntl          ( DownstreamStackBusLane[54][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane25_strm0_data          ( DownstreamStackBusLane[54][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane25_strm0_data_valid    ( DownstreamStackBusLane[54][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane25_strm1_ready         ( DownstreamStackBusLane[54][25].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane25_strm1_cntl          ( DownstreamStackBusLane[54][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane25_strm1_data          ( DownstreamStackBusLane[54][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane25_strm1_data_valid    ( DownstreamStackBusLane[54][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane26_strm0_ready         ( DownstreamStackBusLane[54][26].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane26_strm0_cntl          ( DownstreamStackBusLane[54][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane26_strm0_data          ( DownstreamStackBusLane[54][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane26_strm0_data_valid    ( DownstreamStackBusLane[54][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane26_strm1_ready         ( DownstreamStackBusLane[54][26].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane26_strm1_cntl          ( DownstreamStackBusLane[54][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane26_strm1_data          ( DownstreamStackBusLane[54][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane26_strm1_data_valid    ( DownstreamStackBusLane[54][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane27_strm0_ready         ( DownstreamStackBusLane[54][27].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane27_strm0_cntl          ( DownstreamStackBusLane[54][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane27_strm0_data          ( DownstreamStackBusLane[54][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane27_strm0_data_valid    ( DownstreamStackBusLane[54][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane27_strm1_ready         ( DownstreamStackBusLane[54][27].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane27_strm1_cntl          ( DownstreamStackBusLane[54][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane27_strm1_data          ( DownstreamStackBusLane[54][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane27_strm1_data_valid    ( DownstreamStackBusLane[54][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane28_strm0_ready         ( DownstreamStackBusLane[54][28].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane28_strm0_cntl          ( DownstreamStackBusLane[54][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane28_strm0_data          ( DownstreamStackBusLane[54][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane28_strm0_data_valid    ( DownstreamStackBusLane[54][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane28_strm1_ready         ( DownstreamStackBusLane[54][28].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane28_strm1_cntl          ( DownstreamStackBusLane[54][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane28_strm1_data          ( DownstreamStackBusLane[54][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane28_strm1_data_valid    ( DownstreamStackBusLane[54][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane29_strm0_ready         ( DownstreamStackBusLane[54][29].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane29_strm0_cntl          ( DownstreamStackBusLane[54][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane29_strm0_data          ( DownstreamStackBusLane[54][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane29_strm0_data_valid    ( DownstreamStackBusLane[54][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane29_strm1_ready         ( DownstreamStackBusLane[54][29].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane29_strm1_cntl          ( DownstreamStackBusLane[54][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane29_strm1_data          ( DownstreamStackBusLane[54][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane29_strm1_data_valid    ( DownstreamStackBusLane[54][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane30_strm0_ready         ( DownstreamStackBusLane[54][30].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane30_strm0_cntl          ( DownstreamStackBusLane[54][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane30_strm0_data          ( DownstreamStackBusLane[54][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane30_strm0_data_valid    ( DownstreamStackBusLane[54][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane30_strm1_ready         ( DownstreamStackBusLane[54][30].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane30_strm1_cntl          ( DownstreamStackBusLane[54][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane30_strm1_data          ( DownstreamStackBusLane[54][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane30_strm1_data_valid    ( DownstreamStackBusLane[54][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 54, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane31_strm0_ready         ( DownstreamStackBusLane[54][31].pe__std__lane_strm0_ready              ),      
        .std__pe54__lane31_strm0_cntl          ( DownstreamStackBusLane[54][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe54__lane31_strm0_data          ( DownstreamStackBusLane[54][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe54__lane31_strm0_data_valid    ( DownstreamStackBusLane[54][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__std__lane31_strm1_ready         ( DownstreamStackBusLane[54][31].pe__std__lane_strm1_ready              ),      
        .std__pe54__lane31_strm1_cntl          ( DownstreamStackBusLane[54][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe54__lane31_strm1_data          ( DownstreamStackBusLane[54][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe54__lane31_strm1_data_valid    ( DownstreamStackBusLane[54][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane0_strm0_ready         ( DownstreamStackBusLane[55][0].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane0_strm0_cntl          ( DownstreamStackBusLane[55][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane0_strm0_data          ( DownstreamStackBusLane[55][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane0_strm0_data_valid    ( DownstreamStackBusLane[55][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane0_strm1_ready         ( DownstreamStackBusLane[55][0].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane0_strm1_cntl          ( DownstreamStackBusLane[55][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane0_strm1_data          ( DownstreamStackBusLane[55][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane0_strm1_data_valid    ( DownstreamStackBusLane[55][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane1_strm0_ready         ( DownstreamStackBusLane[55][1].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane1_strm0_cntl          ( DownstreamStackBusLane[55][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane1_strm0_data          ( DownstreamStackBusLane[55][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane1_strm0_data_valid    ( DownstreamStackBusLane[55][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane1_strm1_ready         ( DownstreamStackBusLane[55][1].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane1_strm1_cntl          ( DownstreamStackBusLane[55][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane1_strm1_data          ( DownstreamStackBusLane[55][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane1_strm1_data_valid    ( DownstreamStackBusLane[55][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane2_strm0_ready         ( DownstreamStackBusLane[55][2].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane2_strm0_cntl          ( DownstreamStackBusLane[55][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane2_strm0_data          ( DownstreamStackBusLane[55][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane2_strm0_data_valid    ( DownstreamStackBusLane[55][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane2_strm1_ready         ( DownstreamStackBusLane[55][2].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane2_strm1_cntl          ( DownstreamStackBusLane[55][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane2_strm1_data          ( DownstreamStackBusLane[55][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane2_strm1_data_valid    ( DownstreamStackBusLane[55][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane3_strm0_ready         ( DownstreamStackBusLane[55][3].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane3_strm0_cntl          ( DownstreamStackBusLane[55][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane3_strm0_data          ( DownstreamStackBusLane[55][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane3_strm0_data_valid    ( DownstreamStackBusLane[55][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane3_strm1_ready         ( DownstreamStackBusLane[55][3].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane3_strm1_cntl          ( DownstreamStackBusLane[55][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane3_strm1_data          ( DownstreamStackBusLane[55][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane3_strm1_data_valid    ( DownstreamStackBusLane[55][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane4_strm0_ready         ( DownstreamStackBusLane[55][4].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane4_strm0_cntl          ( DownstreamStackBusLane[55][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane4_strm0_data          ( DownstreamStackBusLane[55][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane4_strm0_data_valid    ( DownstreamStackBusLane[55][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane4_strm1_ready         ( DownstreamStackBusLane[55][4].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane4_strm1_cntl          ( DownstreamStackBusLane[55][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane4_strm1_data          ( DownstreamStackBusLane[55][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane4_strm1_data_valid    ( DownstreamStackBusLane[55][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane5_strm0_ready         ( DownstreamStackBusLane[55][5].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane5_strm0_cntl          ( DownstreamStackBusLane[55][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane5_strm0_data          ( DownstreamStackBusLane[55][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane5_strm0_data_valid    ( DownstreamStackBusLane[55][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane5_strm1_ready         ( DownstreamStackBusLane[55][5].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane5_strm1_cntl          ( DownstreamStackBusLane[55][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane5_strm1_data          ( DownstreamStackBusLane[55][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane5_strm1_data_valid    ( DownstreamStackBusLane[55][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane6_strm0_ready         ( DownstreamStackBusLane[55][6].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane6_strm0_cntl          ( DownstreamStackBusLane[55][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane6_strm0_data          ( DownstreamStackBusLane[55][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane6_strm0_data_valid    ( DownstreamStackBusLane[55][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane6_strm1_ready         ( DownstreamStackBusLane[55][6].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane6_strm1_cntl          ( DownstreamStackBusLane[55][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane6_strm1_data          ( DownstreamStackBusLane[55][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane6_strm1_data_valid    ( DownstreamStackBusLane[55][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane7_strm0_ready         ( DownstreamStackBusLane[55][7].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane7_strm0_cntl          ( DownstreamStackBusLane[55][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane7_strm0_data          ( DownstreamStackBusLane[55][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane7_strm0_data_valid    ( DownstreamStackBusLane[55][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane7_strm1_ready         ( DownstreamStackBusLane[55][7].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane7_strm1_cntl          ( DownstreamStackBusLane[55][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane7_strm1_data          ( DownstreamStackBusLane[55][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane7_strm1_data_valid    ( DownstreamStackBusLane[55][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane8_strm0_ready         ( DownstreamStackBusLane[55][8].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane8_strm0_cntl          ( DownstreamStackBusLane[55][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane8_strm0_data          ( DownstreamStackBusLane[55][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane8_strm0_data_valid    ( DownstreamStackBusLane[55][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane8_strm1_ready         ( DownstreamStackBusLane[55][8].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane8_strm1_cntl          ( DownstreamStackBusLane[55][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane8_strm1_data          ( DownstreamStackBusLane[55][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane8_strm1_data_valid    ( DownstreamStackBusLane[55][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane9_strm0_ready         ( DownstreamStackBusLane[55][9].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane9_strm0_cntl          ( DownstreamStackBusLane[55][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane9_strm0_data          ( DownstreamStackBusLane[55][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane9_strm0_data_valid    ( DownstreamStackBusLane[55][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane9_strm1_ready         ( DownstreamStackBusLane[55][9].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane9_strm1_cntl          ( DownstreamStackBusLane[55][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane9_strm1_data          ( DownstreamStackBusLane[55][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane9_strm1_data_valid    ( DownstreamStackBusLane[55][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane10_strm0_ready         ( DownstreamStackBusLane[55][10].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane10_strm0_cntl          ( DownstreamStackBusLane[55][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane10_strm0_data          ( DownstreamStackBusLane[55][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane10_strm0_data_valid    ( DownstreamStackBusLane[55][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane10_strm1_ready         ( DownstreamStackBusLane[55][10].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane10_strm1_cntl          ( DownstreamStackBusLane[55][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane10_strm1_data          ( DownstreamStackBusLane[55][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane10_strm1_data_valid    ( DownstreamStackBusLane[55][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane11_strm0_ready         ( DownstreamStackBusLane[55][11].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane11_strm0_cntl          ( DownstreamStackBusLane[55][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane11_strm0_data          ( DownstreamStackBusLane[55][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane11_strm0_data_valid    ( DownstreamStackBusLane[55][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane11_strm1_ready         ( DownstreamStackBusLane[55][11].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane11_strm1_cntl          ( DownstreamStackBusLane[55][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane11_strm1_data          ( DownstreamStackBusLane[55][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane11_strm1_data_valid    ( DownstreamStackBusLane[55][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane12_strm0_ready         ( DownstreamStackBusLane[55][12].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane12_strm0_cntl          ( DownstreamStackBusLane[55][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane12_strm0_data          ( DownstreamStackBusLane[55][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane12_strm0_data_valid    ( DownstreamStackBusLane[55][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane12_strm1_ready         ( DownstreamStackBusLane[55][12].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane12_strm1_cntl          ( DownstreamStackBusLane[55][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane12_strm1_data          ( DownstreamStackBusLane[55][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane12_strm1_data_valid    ( DownstreamStackBusLane[55][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane13_strm0_ready         ( DownstreamStackBusLane[55][13].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane13_strm0_cntl          ( DownstreamStackBusLane[55][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane13_strm0_data          ( DownstreamStackBusLane[55][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane13_strm0_data_valid    ( DownstreamStackBusLane[55][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane13_strm1_ready         ( DownstreamStackBusLane[55][13].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane13_strm1_cntl          ( DownstreamStackBusLane[55][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane13_strm1_data          ( DownstreamStackBusLane[55][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane13_strm1_data_valid    ( DownstreamStackBusLane[55][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane14_strm0_ready         ( DownstreamStackBusLane[55][14].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane14_strm0_cntl          ( DownstreamStackBusLane[55][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane14_strm0_data          ( DownstreamStackBusLane[55][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane14_strm0_data_valid    ( DownstreamStackBusLane[55][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane14_strm1_ready         ( DownstreamStackBusLane[55][14].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane14_strm1_cntl          ( DownstreamStackBusLane[55][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane14_strm1_data          ( DownstreamStackBusLane[55][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane14_strm1_data_valid    ( DownstreamStackBusLane[55][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane15_strm0_ready         ( DownstreamStackBusLane[55][15].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane15_strm0_cntl          ( DownstreamStackBusLane[55][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane15_strm0_data          ( DownstreamStackBusLane[55][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane15_strm0_data_valid    ( DownstreamStackBusLane[55][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane15_strm1_ready         ( DownstreamStackBusLane[55][15].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane15_strm1_cntl          ( DownstreamStackBusLane[55][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane15_strm1_data          ( DownstreamStackBusLane[55][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane15_strm1_data_valid    ( DownstreamStackBusLane[55][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane16_strm0_ready         ( DownstreamStackBusLane[55][16].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane16_strm0_cntl          ( DownstreamStackBusLane[55][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane16_strm0_data          ( DownstreamStackBusLane[55][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane16_strm0_data_valid    ( DownstreamStackBusLane[55][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane16_strm1_ready         ( DownstreamStackBusLane[55][16].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane16_strm1_cntl          ( DownstreamStackBusLane[55][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane16_strm1_data          ( DownstreamStackBusLane[55][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane16_strm1_data_valid    ( DownstreamStackBusLane[55][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane17_strm0_ready         ( DownstreamStackBusLane[55][17].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane17_strm0_cntl          ( DownstreamStackBusLane[55][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane17_strm0_data          ( DownstreamStackBusLane[55][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane17_strm0_data_valid    ( DownstreamStackBusLane[55][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane17_strm1_ready         ( DownstreamStackBusLane[55][17].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane17_strm1_cntl          ( DownstreamStackBusLane[55][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane17_strm1_data          ( DownstreamStackBusLane[55][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane17_strm1_data_valid    ( DownstreamStackBusLane[55][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane18_strm0_ready         ( DownstreamStackBusLane[55][18].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane18_strm0_cntl          ( DownstreamStackBusLane[55][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane18_strm0_data          ( DownstreamStackBusLane[55][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane18_strm0_data_valid    ( DownstreamStackBusLane[55][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane18_strm1_ready         ( DownstreamStackBusLane[55][18].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane18_strm1_cntl          ( DownstreamStackBusLane[55][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane18_strm1_data          ( DownstreamStackBusLane[55][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane18_strm1_data_valid    ( DownstreamStackBusLane[55][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane19_strm0_ready         ( DownstreamStackBusLane[55][19].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane19_strm0_cntl          ( DownstreamStackBusLane[55][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane19_strm0_data          ( DownstreamStackBusLane[55][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane19_strm0_data_valid    ( DownstreamStackBusLane[55][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane19_strm1_ready         ( DownstreamStackBusLane[55][19].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane19_strm1_cntl          ( DownstreamStackBusLane[55][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane19_strm1_data          ( DownstreamStackBusLane[55][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane19_strm1_data_valid    ( DownstreamStackBusLane[55][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane20_strm0_ready         ( DownstreamStackBusLane[55][20].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane20_strm0_cntl          ( DownstreamStackBusLane[55][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane20_strm0_data          ( DownstreamStackBusLane[55][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane20_strm0_data_valid    ( DownstreamStackBusLane[55][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane20_strm1_ready         ( DownstreamStackBusLane[55][20].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane20_strm1_cntl          ( DownstreamStackBusLane[55][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane20_strm1_data          ( DownstreamStackBusLane[55][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane20_strm1_data_valid    ( DownstreamStackBusLane[55][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane21_strm0_ready         ( DownstreamStackBusLane[55][21].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane21_strm0_cntl          ( DownstreamStackBusLane[55][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane21_strm0_data          ( DownstreamStackBusLane[55][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane21_strm0_data_valid    ( DownstreamStackBusLane[55][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane21_strm1_ready         ( DownstreamStackBusLane[55][21].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane21_strm1_cntl          ( DownstreamStackBusLane[55][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane21_strm1_data          ( DownstreamStackBusLane[55][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane21_strm1_data_valid    ( DownstreamStackBusLane[55][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane22_strm0_ready         ( DownstreamStackBusLane[55][22].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane22_strm0_cntl          ( DownstreamStackBusLane[55][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane22_strm0_data          ( DownstreamStackBusLane[55][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane22_strm0_data_valid    ( DownstreamStackBusLane[55][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane22_strm1_ready         ( DownstreamStackBusLane[55][22].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane22_strm1_cntl          ( DownstreamStackBusLane[55][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane22_strm1_data          ( DownstreamStackBusLane[55][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane22_strm1_data_valid    ( DownstreamStackBusLane[55][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane23_strm0_ready         ( DownstreamStackBusLane[55][23].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane23_strm0_cntl          ( DownstreamStackBusLane[55][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane23_strm0_data          ( DownstreamStackBusLane[55][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane23_strm0_data_valid    ( DownstreamStackBusLane[55][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane23_strm1_ready         ( DownstreamStackBusLane[55][23].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane23_strm1_cntl          ( DownstreamStackBusLane[55][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane23_strm1_data          ( DownstreamStackBusLane[55][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane23_strm1_data_valid    ( DownstreamStackBusLane[55][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane24_strm0_ready         ( DownstreamStackBusLane[55][24].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane24_strm0_cntl          ( DownstreamStackBusLane[55][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane24_strm0_data          ( DownstreamStackBusLane[55][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane24_strm0_data_valid    ( DownstreamStackBusLane[55][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane24_strm1_ready         ( DownstreamStackBusLane[55][24].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane24_strm1_cntl          ( DownstreamStackBusLane[55][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane24_strm1_data          ( DownstreamStackBusLane[55][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane24_strm1_data_valid    ( DownstreamStackBusLane[55][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane25_strm0_ready         ( DownstreamStackBusLane[55][25].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane25_strm0_cntl          ( DownstreamStackBusLane[55][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane25_strm0_data          ( DownstreamStackBusLane[55][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane25_strm0_data_valid    ( DownstreamStackBusLane[55][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane25_strm1_ready         ( DownstreamStackBusLane[55][25].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane25_strm1_cntl          ( DownstreamStackBusLane[55][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane25_strm1_data          ( DownstreamStackBusLane[55][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane25_strm1_data_valid    ( DownstreamStackBusLane[55][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane26_strm0_ready         ( DownstreamStackBusLane[55][26].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane26_strm0_cntl          ( DownstreamStackBusLane[55][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane26_strm0_data          ( DownstreamStackBusLane[55][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane26_strm0_data_valid    ( DownstreamStackBusLane[55][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane26_strm1_ready         ( DownstreamStackBusLane[55][26].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane26_strm1_cntl          ( DownstreamStackBusLane[55][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane26_strm1_data          ( DownstreamStackBusLane[55][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane26_strm1_data_valid    ( DownstreamStackBusLane[55][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane27_strm0_ready         ( DownstreamStackBusLane[55][27].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane27_strm0_cntl          ( DownstreamStackBusLane[55][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane27_strm0_data          ( DownstreamStackBusLane[55][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane27_strm0_data_valid    ( DownstreamStackBusLane[55][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane27_strm1_ready         ( DownstreamStackBusLane[55][27].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane27_strm1_cntl          ( DownstreamStackBusLane[55][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane27_strm1_data          ( DownstreamStackBusLane[55][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane27_strm1_data_valid    ( DownstreamStackBusLane[55][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane28_strm0_ready         ( DownstreamStackBusLane[55][28].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane28_strm0_cntl          ( DownstreamStackBusLane[55][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane28_strm0_data          ( DownstreamStackBusLane[55][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane28_strm0_data_valid    ( DownstreamStackBusLane[55][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane28_strm1_ready         ( DownstreamStackBusLane[55][28].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane28_strm1_cntl          ( DownstreamStackBusLane[55][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane28_strm1_data          ( DownstreamStackBusLane[55][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane28_strm1_data_valid    ( DownstreamStackBusLane[55][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane29_strm0_ready         ( DownstreamStackBusLane[55][29].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane29_strm0_cntl          ( DownstreamStackBusLane[55][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane29_strm0_data          ( DownstreamStackBusLane[55][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane29_strm0_data_valid    ( DownstreamStackBusLane[55][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane29_strm1_ready         ( DownstreamStackBusLane[55][29].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane29_strm1_cntl          ( DownstreamStackBusLane[55][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane29_strm1_data          ( DownstreamStackBusLane[55][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane29_strm1_data_valid    ( DownstreamStackBusLane[55][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane30_strm0_ready         ( DownstreamStackBusLane[55][30].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane30_strm0_cntl          ( DownstreamStackBusLane[55][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane30_strm0_data          ( DownstreamStackBusLane[55][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane30_strm0_data_valid    ( DownstreamStackBusLane[55][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane30_strm1_ready         ( DownstreamStackBusLane[55][30].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane30_strm1_cntl          ( DownstreamStackBusLane[55][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane30_strm1_data          ( DownstreamStackBusLane[55][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane30_strm1_data_valid    ( DownstreamStackBusLane[55][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 55, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane31_strm0_ready         ( DownstreamStackBusLane[55][31].pe__std__lane_strm0_ready              ),      
        .std__pe55__lane31_strm0_cntl          ( DownstreamStackBusLane[55][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe55__lane31_strm0_data          ( DownstreamStackBusLane[55][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe55__lane31_strm0_data_valid    ( DownstreamStackBusLane[55][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__std__lane31_strm1_ready         ( DownstreamStackBusLane[55][31].pe__std__lane_strm1_ready              ),      
        .std__pe55__lane31_strm1_cntl          ( DownstreamStackBusLane[55][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe55__lane31_strm1_data          ( DownstreamStackBusLane[55][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe55__lane31_strm1_data_valid    ( DownstreamStackBusLane[55][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane0_strm0_ready         ( DownstreamStackBusLane[56][0].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane0_strm0_cntl          ( DownstreamStackBusLane[56][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane0_strm0_data          ( DownstreamStackBusLane[56][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane0_strm0_data_valid    ( DownstreamStackBusLane[56][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane0_strm1_ready         ( DownstreamStackBusLane[56][0].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane0_strm1_cntl          ( DownstreamStackBusLane[56][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane0_strm1_data          ( DownstreamStackBusLane[56][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane0_strm1_data_valid    ( DownstreamStackBusLane[56][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane1_strm0_ready         ( DownstreamStackBusLane[56][1].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane1_strm0_cntl          ( DownstreamStackBusLane[56][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane1_strm0_data          ( DownstreamStackBusLane[56][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane1_strm0_data_valid    ( DownstreamStackBusLane[56][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane1_strm1_ready         ( DownstreamStackBusLane[56][1].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane1_strm1_cntl          ( DownstreamStackBusLane[56][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane1_strm1_data          ( DownstreamStackBusLane[56][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane1_strm1_data_valid    ( DownstreamStackBusLane[56][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane2_strm0_ready         ( DownstreamStackBusLane[56][2].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane2_strm0_cntl          ( DownstreamStackBusLane[56][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane2_strm0_data          ( DownstreamStackBusLane[56][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane2_strm0_data_valid    ( DownstreamStackBusLane[56][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane2_strm1_ready         ( DownstreamStackBusLane[56][2].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane2_strm1_cntl          ( DownstreamStackBusLane[56][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane2_strm1_data          ( DownstreamStackBusLane[56][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane2_strm1_data_valid    ( DownstreamStackBusLane[56][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane3_strm0_ready         ( DownstreamStackBusLane[56][3].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane3_strm0_cntl          ( DownstreamStackBusLane[56][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane3_strm0_data          ( DownstreamStackBusLane[56][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane3_strm0_data_valid    ( DownstreamStackBusLane[56][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane3_strm1_ready         ( DownstreamStackBusLane[56][3].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane3_strm1_cntl          ( DownstreamStackBusLane[56][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane3_strm1_data          ( DownstreamStackBusLane[56][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane3_strm1_data_valid    ( DownstreamStackBusLane[56][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane4_strm0_ready         ( DownstreamStackBusLane[56][4].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane4_strm0_cntl          ( DownstreamStackBusLane[56][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane4_strm0_data          ( DownstreamStackBusLane[56][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane4_strm0_data_valid    ( DownstreamStackBusLane[56][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane4_strm1_ready         ( DownstreamStackBusLane[56][4].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane4_strm1_cntl          ( DownstreamStackBusLane[56][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane4_strm1_data          ( DownstreamStackBusLane[56][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane4_strm1_data_valid    ( DownstreamStackBusLane[56][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane5_strm0_ready         ( DownstreamStackBusLane[56][5].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane5_strm0_cntl          ( DownstreamStackBusLane[56][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane5_strm0_data          ( DownstreamStackBusLane[56][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane5_strm0_data_valid    ( DownstreamStackBusLane[56][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane5_strm1_ready         ( DownstreamStackBusLane[56][5].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane5_strm1_cntl          ( DownstreamStackBusLane[56][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane5_strm1_data          ( DownstreamStackBusLane[56][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane5_strm1_data_valid    ( DownstreamStackBusLane[56][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane6_strm0_ready         ( DownstreamStackBusLane[56][6].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane6_strm0_cntl          ( DownstreamStackBusLane[56][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane6_strm0_data          ( DownstreamStackBusLane[56][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane6_strm0_data_valid    ( DownstreamStackBusLane[56][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane6_strm1_ready         ( DownstreamStackBusLane[56][6].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane6_strm1_cntl          ( DownstreamStackBusLane[56][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane6_strm1_data          ( DownstreamStackBusLane[56][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane6_strm1_data_valid    ( DownstreamStackBusLane[56][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane7_strm0_ready         ( DownstreamStackBusLane[56][7].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane7_strm0_cntl          ( DownstreamStackBusLane[56][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane7_strm0_data          ( DownstreamStackBusLane[56][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane7_strm0_data_valid    ( DownstreamStackBusLane[56][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane7_strm1_ready         ( DownstreamStackBusLane[56][7].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane7_strm1_cntl          ( DownstreamStackBusLane[56][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane7_strm1_data          ( DownstreamStackBusLane[56][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane7_strm1_data_valid    ( DownstreamStackBusLane[56][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane8_strm0_ready         ( DownstreamStackBusLane[56][8].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane8_strm0_cntl          ( DownstreamStackBusLane[56][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane8_strm0_data          ( DownstreamStackBusLane[56][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane8_strm0_data_valid    ( DownstreamStackBusLane[56][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane8_strm1_ready         ( DownstreamStackBusLane[56][8].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane8_strm1_cntl          ( DownstreamStackBusLane[56][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane8_strm1_data          ( DownstreamStackBusLane[56][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane8_strm1_data_valid    ( DownstreamStackBusLane[56][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane9_strm0_ready         ( DownstreamStackBusLane[56][9].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane9_strm0_cntl          ( DownstreamStackBusLane[56][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane9_strm0_data          ( DownstreamStackBusLane[56][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane9_strm0_data_valid    ( DownstreamStackBusLane[56][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane9_strm1_ready         ( DownstreamStackBusLane[56][9].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane9_strm1_cntl          ( DownstreamStackBusLane[56][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane9_strm1_data          ( DownstreamStackBusLane[56][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane9_strm1_data_valid    ( DownstreamStackBusLane[56][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane10_strm0_ready         ( DownstreamStackBusLane[56][10].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane10_strm0_cntl          ( DownstreamStackBusLane[56][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane10_strm0_data          ( DownstreamStackBusLane[56][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane10_strm0_data_valid    ( DownstreamStackBusLane[56][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane10_strm1_ready         ( DownstreamStackBusLane[56][10].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane10_strm1_cntl          ( DownstreamStackBusLane[56][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane10_strm1_data          ( DownstreamStackBusLane[56][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane10_strm1_data_valid    ( DownstreamStackBusLane[56][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane11_strm0_ready         ( DownstreamStackBusLane[56][11].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane11_strm0_cntl          ( DownstreamStackBusLane[56][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane11_strm0_data          ( DownstreamStackBusLane[56][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane11_strm0_data_valid    ( DownstreamStackBusLane[56][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane11_strm1_ready         ( DownstreamStackBusLane[56][11].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane11_strm1_cntl          ( DownstreamStackBusLane[56][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane11_strm1_data          ( DownstreamStackBusLane[56][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane11_strm1_data_valid    ( DownstreamStackBusLane[56][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane12_strm0_ready         ( DownstreamStackBusLane[56][12].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane12_strm0_cntl          ( DownstreamStackBusLane[56][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane12_strm0_data          ( DownstreamStackBusLane[56][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane12_strm0_data_valid    ( DownstreamStackBusLane[56][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane12_strm1_ready         ( DownstreamStackBusLane[56][12].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane12_strm1_cntl          ( DownstreamStackBusLane[56][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane12_strm1_data          ( DownstreamStackBusLane[56][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane12_strm1_data_valid    ( DownstreamStackBusLane[56][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane13_strm0_ready         ( DownstreamStackBusLane[56][13].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane13_strm0_cntl          ( DownstreamStackBusLane[56][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane13_strm0_data          ( DownstreamStackBusLane[56][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane13_strm0_data_valid    ( DownstreamStackBusLane[56][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane13_strm1_ready         ( DownstreamStackBusLane[56][13].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane13_strm1_cntl          ( DownstreamStackBusLane[56][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane13_strm1_data          ( DownstreamStackBusLane[56][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane13_strm1_data_valid    ( DownstreamStackBusLane[56][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane14_strm0_ready         ( DownstreamStackBusLane[56][14].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane14_strm0_cntl          ( DownstreamStackBusLane[56][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane14_strm0_data          ( DownstreamStackBusLane[56][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane14_strm0_data_valid    ( DownstreamStackBusLane[56][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane14_strm1_ready         ( DownstreamStackBusLane[56][14].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane14_strm1_cntl          ( DownstreamStackBusLane[56][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane14_strm1_data          ( DownstreamStackBusLane[56][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane14_strm1_data_valid    ( DownstreamStackBusLane[56][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane15_strm0_ready         ( DownstreamStackBusLane[56][15].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane15_strm0_cntl          ( DownstreamStackBusLane[56][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane15_strm0_data          ( DownstreamStackBusLane[56][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane15_strm0_data_valid    ( DownstreamStackBusLane[56][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane15_strm1_ready         ( DownstreamStackBusLane[56][15].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane15_strm1_cntl          ( DownstreamStackBusLane[56][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane15_strm1_data          ( DownstreamStackBusLane[56][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane15_strm1_data_valid    ( DownstreamStackBusLane[56][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane16_strm0_ready         ( DownstreamStackBusLane[56][16].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane16_strm0_cntl          ( DownstreamStackBusLane[56][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane16_strm0_data          ( DownstreamStackBusLane[56][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane16_strm0_data_valid    ( DownstreamStackBusLane[56][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane16_strm1_ready         ( DownstreamStackBusLane[56][16].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane16_strm1_cntl          ( DownstreamStackBusLane[56][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane16_strm1_data          ( DownstreamStackBusLane[56][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane16_strm1_data_valid    ( DownstreamStackBusLane[56][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane17_strm0_ready         ( DownstreamStackBusLane[56][17].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane17_strm0_cntl          ( DownstreamStackBusLane[56][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane17_strm0_data          ( DownstreamStackBusLane[56][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane17_strm0_data_valid    ( DownstreamStackBusLane[56][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane17_strm1_ready         ( DownstreamStackBusLane[56][17].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane17_strm1_cntl          ( DownstreamStackBusLane[56][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane17_strm1_data          ( DownstreamStackBusLane[56][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane17_strm1_data_valid    ( DownstreamStackBusLane[56][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane18_strm0_ready         ( DownstreamStackBusLane[56][18].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane18_strm0_cntl          ( DownstreamStackBusLane[56][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane18_strm0_data          ( DownstreamStackBusLane[56][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane18_strm0_data_valid    ( DownstreamStackBusLane[56][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane18_strm1_ready         ( DownstreamStackBusLane[56][18].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane18_strm1_cntl          ( DownstreamStackBusLane[56][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane18_strm1_data          ( DownstreamStackBusLane[56][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane18_strm1_data_valid    ( DownstreamStackBusLane[56][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane19_strm0_ready         ( DownstreamStackBusLane[56][19].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane19_strm0_cntl          ( DownstreamStackBusLane[56][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane19_strm0_data          ( DownstreamStackBusLane[56][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane19_strm0_data_valid    ( DownstreamStackBusLane[56][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane19_strm1_ready         ( DownstreamStackBusLane[56][19].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane19_strm1_cntl          ( DownstreamStackBusLane[56][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane19_strm1_data          ( DownstreamStackBusLane[56][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane19_strm1_data_valid    ( DownstreamStackBusLane[56][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane20_strm0_ready         ( DownstreamStackBusLane[56][20].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane20_strm0_cntl          ( DownstreamStackBusLane[56][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane20_strm0_data          ( DownstreamStackBusLane[56][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane20_strm0_data_valid    ( DownstreamStackBusLane[56][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane20_strm1_ready         ( DownstreamStackBusLane[56][20].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane20_strm1_cntl          ( DownstreamStackBusLane[56][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane20_strm1_data          ( DownstreamStackBusLane[56][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane20_strm1_data_valid    ( DownstreamStackBusLane[56][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane21_strm0_ready         ( DownstreamStackBusLane[56][21].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane21_strm0_cntl          ( DownstreamStackBusLane[56][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane21_strm0_data          ( DownstreamStackBusLane[56][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane21_strm0_data_valid    ( DownstreamStackBusLane[56][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane21_strm1_ready         ( DownstreamStackBusLane[56][21].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane21_strm1_cntl          ( DownstreamStackBusLane[56][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane21_strm1_data          ( DownstreamStackBusLane[56][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane21_strm1_data_valid    ( DownstreamStackBusLane[56][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane22_strm0_ready         ( DownstreamStackBusLane[56][22].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane22_strm0_cntl          ( DownstreamStackBusLane[56][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane22_strm0_data          ( DownstreamStackBusLane[56][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane22_strm0_data_valid    ( DownstreamStackBusLane[56][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane22_strm1_ready         ( DownstreamStackBusLane[56][22].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane22_strm1_cntl          ( DownstreamStackBusLane[56][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane22_strm1_data          ( DownstreamStackBusLane[56][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane22_strm1_data_valid    ( DownstreamStackBusLane[56][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane23_strm0_ready         ( DownstreamStackBusLane[56][23].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane23_strm0_cntl          ( DownstreamStackBusLane[56][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane23_strm0_data          ( DownstreamStackBusLane[56][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane23_strm0_data_valid    ( DownstreamStackBusLane[56][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane23_strm1_ready         ( DownstreamStackBusLane[56][23].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane23_strm1_cntl          ( DownstreamStackBusLane[56][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane23_strm1_data          ( DownstreamStackBusLane[56][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane23_strm1_data_valid    ( DownstreamStackBusLane[56][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane24_strm0_ready         ( DownstreamStackBusLane[56][24].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane24_strm0_cntl          ( DownstreamStackBusLane[56][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane24_strm0_data          ( DownstreamStackBusLane[56][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane24_strm0_data_valid    ( DownstreamStackBusLane[56][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane24_strm1_ready         ( DownstreamStackBusLane[56][24].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane24_strm1_cntl          ( DownstreamStackBusLane[56][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane24_strm1_data          ( DownstreamStackBusLane[56][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane24_strm1_data_valid    ( DownstreamStackBusLane[56][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane25_strm0_ready         ( DownstreamStackBusLane[56][25].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane25_strm0_cntl          ( DownstreamStackBusLane[56][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane25_strm0_data          ( DownstreamStackBusLane[56][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane25_strm0_data_valid    ( DownstreamStackBusLane[56][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane25_strm1_ready         ( DownstreamStackBusLane[56][25].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane25_strm1_cntl          ( DownstreamStackBusLane[56][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane25_strm1_data          ( DownstreamStackBusLane[56][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane25_strm1_data_valid    ( DownstreamStackBusLane[56][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane26_strm0_ready         ( DownstreamStackBusLane[56][26].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane26_strm0_cntl          ( DownstreamStackBusLane[56][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane26_strm0_data          ( DownstreamStackBusLane[56][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane26_strm0_data_valid    ( DownstreamStackBusLane[56][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane26_strm1_ready         ( DownstreamStackBusLane[56][26].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane26_strm1_cntl          ( DownstreamStackBusLane[56][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane26_strm1_data          ( DownstreamStackBusLane[56][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane26_strm1_data_valid    ( DownstreamStackBusLane[56][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane27_strm0_ready         ( DownstreamStackBusLane[56][27].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane27_strm0_cntl          ( DownstreamStackBusLane[56][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane27_strm0_data          ( DownstreamStackBusLane[56][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane27_strm0_data_valid    ( DownstreamStackBusLane[56][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane27_strm1_ready         ( DownstreamStackBusLane[56][27].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane27_strm1_cntl          ( DownstreamStackBusLane[56][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane27_strm1_data          ( DownstreamStackBusLane[56][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane27_strm1_data_valid    ( DownstreamStackBusLane[56][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane28_strm0_ready         ( DownstreamStackBusLane[56][28].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane28_strm0_cntl          ( DownstreamStackBusLane[56][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane28_strm0_data          ( DownstreamStackBusLane[56][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane28_strm0_data_valid    ( DownstreamStackBusLane[56][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane28_strm1_ready         ( DownstreamStackBusLane[56][28].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane28_strm1_cntl          ( DownstreamStackBusLane[56][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane28_strm1_data          ( DownstreamStackBusLane[56][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane28_strm1_data_valid    ( DownstreamStackBusLane[56][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane29_strm0_ready         ( DownstreamStackBusLane[56][29].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane29_strm0_cntl          ( DownstreamStackBusLane[56][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane29_strm0_data          ( DownstreamStackBusLane[56][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane29_strm0_data_valid    ( DownstreamStackBusLane[56][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane29_strm1_ready         ( DownstreamStackBusLane[56][29].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane29_strm1_cntl          ( DownstreamStackBusLane[56][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane29_strm1_data          ( DownstreamStackBusLane[56][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane29_strm1_data_valid    ( DownstreamStackBusLane[56][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane30_strm0_ready         ( DownstreamStackBusLane[56][30].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane30_strm0_cntl          ( DownstreamStackBusLane[56][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane30_strm0_data          ( DownstreamStackBusLane[56][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane30_strm0_data_valid    ( DownstreamStackBusLane[56][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane30_strm1_ready         ( DownstreamStackBusLane[56][30].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane30_strm1_cntl          ( DownstreamStackBusLane[56][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane30_strm1_data          ( DownstreamStackBusLane[56][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane30_strm1_data_valid    ( DownstreamStackBusLane[56][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 56, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane31_strm0_ready         ( DownstreamStackBusLane[56][31].pe__std__lane_strm0_ready              ),      
        .std__pe56__lane31_strm0_cntl          ( DownstreamStackBusLane[56][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe56__lane31_strm0_data          ( DownstreamStackBusLane[56][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe56__lane31_strm0_data_valid    ( DownstreamStackBusLane[56][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__std__lane31_strm1_ready         ( DownstreamStackBusLane[56][31].pe__std__lane_strm1_ready              ),      
        .std__pe56__lane31_strm1_cntl          ( DownstreamStackBusLane[56][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe56__lane31_strm1_data          ( DownstreamStackBusLane[56][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe56__lane31_strm1_data_valid    ( DownstreamStackBusLane[56][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane0_strm0_ready         ( DownstreamStackBusLane[57][0].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane0_strm0_cntl          ( DownstreamStackBusLane[57][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane0_strm0_data          ( DownstreamStackBusLane[57][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane0_strm0_data_valid    ( DownstreamStackBusLane[57][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane0_strm1_ready         ( DownstreamStackBusLane[57][0].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane0_strm1_cntl          ( DownstreamStackBusLane[57][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane0_strm1_data          ( DownstreamStackBusLane[57][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane0_strm1_data_valid    ( DownstreamStackBusLane[57][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane1_strm0_ready         ( DownstreamStackBusLane[57][1].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane1_strm0_cntl          ( DownstreamStackBusLane[57][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane1_strm0_data          ( DownstreamStackBusLane[57][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane1_strm0_data_valid    ( DownstreamStackBusLane[57][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane1_strm1_ready         ( DownstreamStackBusLane[57][1].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane1_strm1_cntl          ( DownstreamStackBusLane[57][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane1_strm1_data          ( DownstreamStackBusLane[57][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane1_strm1_data_valid    ( DownstreamStackBusLane[57][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane2_strm0_ready         ( DownstreamStackBusLane[57][2].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane2_strm0_cntl          ( DownstreamStackBusLane[57][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane2_strm0_data          ( DownstreamStackBusLane[57][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane2_strm0_data_valid    ( DownstreamStackBusLane[57][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane2_strm1_ready         ( DownstreamStackBusLane[57][2].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane2_strm1_cntl          ( DownstreamStackBusLane[57][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane2_strm1_data          ( DownstreamStackBusLane[57][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane2_strm1_data_valid    ( DownstreamStackBusLane[57][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane3_strm0_ready         ( DownstreamStackBusLane[57][3].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane3_strm0_cntl          ( DownstreamStackBusLane[57][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane3_strm0_data          ( DownstreamStackBusLane[57][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane3_strm0_data_valid    ( DownstreamStackBusLane[57][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane3_strm1_ready         ( DownstreamStackBusLane[57][3].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane3_strm1_cntl          ( DownstreamStackBusLane[57][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane3_strm1_data          ( DownstreamStackBusLane[57][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane3_strm1_data_valid    ( DownstreamStackBusLane[57][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane4_strm0_ready         ( DownstreamStackBusLane[57][4].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane4_strm0_cntl          ( DownstreamStackBusLane[57][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane4_strm0_data          ( DownstreamStackBusLane[57][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane4_strm0_data_valid    ( DownstreamStackBusLane[57][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane4_strm1_ready         ( DownstreamStackBusLane[57][4].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane4_strm1_cntl          ( DownstreamStackBusLane[57][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane4_strm1_data          ( DownstreamStackBusLane[57][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane4_strm1_data_valid    ( DownstreamStackBusLane[57][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane5_strm0_ready         ( DownstreamStackBusLane[57][5].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane5_strm0_cntl          ( DownstreamStackBusLane[57][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane5_strm0_data          ( DownstreamStackBusLane[57][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane5_strm0_data_valid    ( DownstreamStackBusLane[57][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane5_strm1_ready         ( DownstreamStackBusLane[57][5].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane5_strm1_cntl          ( DownstreamStackBusLane[57][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane5_strm1_data          ( DownstreamStackBusLane[57][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane5_strm1_data_valid    ( DownstreamStackBusLane[57][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane6_strm0_ready         ( DownstreamStackBusLane[57][6].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane6_strm0_cntl          ( DownstreamStackBusLane[57][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane6_strm0_data          ( DownstreamStackBusLane[57][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane6_strm0_data_valid    ( DownstreamStackBusLane[57][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane6_strm1_ready         ( DownstreamStackBusLane[57][6].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane6_strm1_cntl          ( DownstreamStackBusLane[57][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane6_strm1_data          ( DownstreamStackBusLane[57][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane6_strm1_data_valid    ( DownstreamStackBusLane[57][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane7_strm0_ready         ( DownstreamStackBusLane[57][7].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane7_strm0_cntl          ( DownstreamStackBusLane[57][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane7_strm0_data          ( DownstreamStackBusLane[57][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane7_strm0_data_valid    ( DownstreamStackBusLane[57][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane7_strm1_ready         ( DownstreamStackBusLane[57][7].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane7_strm1_cntl          ( DownstreamStackBusLane[57][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane7_strm1_data          ( DownstreamStackBusLane[57][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane7_strm1_data_valid    ( DownstreamStackBusLane[57][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane8_strm0_ready         ( DownstreamStackBusLane[57][8].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane8_strm0_cntl          ( DownstreamStackBusLane[57][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane8_strm0_data          ( DownstreamStackBusLane[57][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane8_strm0_data_valid    ( DownstreamStackBusLane[57][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane8_strm1_ready         ( DownstreamStackBusLane[57][8].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane8_strm1_cntl          ( DownstreamStackBusLane[57][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane8_strm1_data          ( DownstreamStackBusLane[57][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane8_strm1_data_valid    ( DownstreamStackBusLane[57][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane9_strm0_ready         ( DownstreamStackBusLane[57][9].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane9_strm0_cntl          ( DownstreamStackBusLane[57][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane9_strm0_data          ( DownstreamStackBusLane[57][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane9_strm0_data_valid    ( DownstreamStackBusLane[57][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane9_strm1_ready         ( DownstreamStackBusLane[57][9].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane9_strm1_cntl          ( DownstreamStackBusLane[57][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane9_strm1_data          ( DownstreamStackBusLane[57][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane9_strm1_data_valid    ( DownstreamStackBusLane[57][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane10_strm0_ready         ( DownstreamStackBusLane[57][10].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane10_strm0_cntl          ( DownstreamStackBusLane[57][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane10_strm0_data          ( DownstreamStackBusLane[57][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane10_strm0_data_valid    ( DownstreamStackBusLane[57][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane10_strm1_ready         ( DownstreamStackBusLane[57][10].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane10_strm1_cntl          ( DownstreamStackBusLane[57][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane10_strm1_data          ( DownstreamStackBusLane[57][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane10_strm1_data_valid    ( DownstreamStackBusLane[57][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane11_strm0_ready         ( DownstreamStackBusLane[57][11].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane11_strm0_cntl          ( DownstreamStackBusLane[57][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane11_strm0_data          ( DownstreamStackBusLane[57][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane11_strm0_data_valid    ( DownstreamStackBusLane[57][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane11_strm1_ready         ( DownstreamStackBusLane[57][11].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane11_strm1_cntl          ( DownstreamStackBusLane[57][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane11_strm1_data          ( DownstreamStackBusLane[57][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane11_strm1_data_valid    ( DownstreamStackBusLane[57][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane12_strm0_ready         ( DownstreamStackBusLane[57][12].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane12_strm0_cntl          ( DownstreamStackBusLane[57][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane12_strm0_data          ( DownstreamStackBusLane[57][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane12_strm0_data_valid    ( DownstreamStackBusLane[57][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane12_strm1_ready         ( DownstreamStackBusLane[57][12].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane12_strm1_cntl          ( DownstreamStackBusLane[57][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane12_strm1_data          ( DownstreamStackBusLane[57][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane12_strm1_data_valid    ( DownstreamStackBusLane[57][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane13_strm0_ready         ( DownstreamStackBusLane[57][13].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane13_strm0_cntl          ( DownstreamStackBusLane[57][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane13_strm0_data          ( DownstreamStackBusLane[57][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane13_strm0_data_valid    ( DownstreamStackBusLane[57][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane13_strm1_ready         ( DownstreamStackBusLane[57][13].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane13_strm1_cntl          ( DownstreamStackBusLane[57][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane13_strm1_data          ( DownstreamStackBusLane[57][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane13_strm1_data_valid    ( DownstreamStackBusLane[57][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane14_strm0_ready         ( DownstreamStackBusLane[57][14].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane14_strm0_cntl          ( DownstreamStackBusLane[57][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane14_strm0_data          ( DownstreamStackBusLane[57][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane14_strm0_data_valid    ( DownstreamStackBusLane[57][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane14_strm1_ready         ( DownstreamStackBusLane[57][14].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane14_strm1_cntl          ( DownstreamStackBusLane[57][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane14_strm1_data          ( DownstreamStackBusLane[57][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane14_strm1_data_valid    ( DownstreamStackBusLane[57][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane15_strm0_ready         ( DownstreamStackBusLane[57][15].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane15_strm0_cntl          ( DownstreamStackBusLane[57][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane15_strm0_data          ( DownstreamStackBusLane[57][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane15_strm0_data_valid    ( DownstreamStackBusLane[57][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane15_strm1_ready         ( DownstreamStackBusLane[57][15].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane15_strm1_cntl          ( DownstreamStackBusLane[57][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane15_strm1_data          ( DownstreamStackBusLane[57][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane15_strm1_data_valid    ( DownstreamStackBusLane[57][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane16_strm0_ready         ( DownstreamStackBusLane[57][16].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane16_strm0_cntl          ( DownstreamStackBusLane[57][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane16_strm0_data          ( DownstreamStackBusLane[57][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane16_strm0_data_valid    ( DownstreamStackBusLane[57][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane16_strm1_ready         ( DownstreamStackBusLane[57][16].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane16_strm1_cntl          ( DownstreamStackBusLane[57][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane16_strm1_data          ( DownstreamStackBusLane[57][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane16_strm1_data_valid    ( DownstreamStackBusLane[57][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane17_strm0_ready         ( DownstreamStackBusLane[57][17].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane17_strm0_cntl          ( DownstreamStackBusLane[57][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane17_strm0_data          ( DownstreamStackBusLane[57][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane17_strm0_data_valid    ( DownstreamStackBusLane[57][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane17_strm1_ready         ( DownstreamStackBusLane[57][17].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane17_strm1_cntl          ( DownstreamStackBusLane[57][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane17_strm1_data          ( DownstreamStackBusLane[57][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane17_strm1_data_valid    ( DownstreamStackBusLane[57][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane18_strm0_ready         ( DownstreamStackBusLane[57][18].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane18_strm0_cntl          ( DownstreamStackBusLane[57][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane18_strm0_data          ( DownstreamStackBusLane[57][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane18_strm0_data_valid    ( DownstreamStackBusLane[57][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane18_strm1_ready         ( DownstreamStackBusLane[57][18].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane18_strm1_cntl          ( DownstreamStackBusLane[57][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane18_strm1_data          ( DownstreamStackBusLane[57][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane18_strm1_data_valid    ( DownstreamStackBusLane[57][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane19_strm0_ready         ( DownstreamStackBusLane[57][19].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane19_strm0_cntl          ( DownstreamStackBusLane[57][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane19_strm0_data          ( DownstreamStackBusLane[57][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane19_strm0_data_valid    ( DownstreamStackBusLane[57][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane19_strm1_ready         ( DownstreamStackBusLane[57][19].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane19_strm1_cntl          ( DownstreamStackBusLane[57][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane19_strm1_data          ( DownstreamStackBusLane[57][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane19_strm1_data_valid    ( DownstreamStackBusLane[57][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane20_strm0_ready         ( DownstreamStackBusLane[57][20].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane20_strm0_cntl          ( DownstreamStackBusLane[57][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane20_strm0_data          ( DownstreamStackBusLane[57][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane20_strm0_data_valid    ( DownstreamStackBusLane[57][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane20_strm1_ready         ( DownstreamStackBusLane[57][20].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane20_strm1_cntl          ( DownstreamStackBusLane[57][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane20_strm1_data          ( DownstreamStackBusLane[57][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane20_strm1_data_valid    ( DownstreamStackBusLane[57][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane21_strm0_ready         ( DownstreamStackBusLane[57][21].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane21_strm0_cntl          ( DownstreamStackBusLane[57][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane21_strm0_data          ( DownstreamStackBusLane[57][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane21_strm0_data_valid    ( DownstreamStackBusLane[57][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane21_strm1_ready         ( DownstreamStackBusLane[57][21].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane21_strm1_cntl          ( DownstreamStackBusLane[57][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane21_strm1_data          ( DownstreamStackBusLane[57][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane21_strm1_data_valid    ( DownstreamStackBusLane[57][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane22_strm0_ready         ( DownstreamStackBusLane[57][22].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane22_strm0_cntl          ( DownstreamStackBusLane[57][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane22_strm0_data          ( DownstreamStackBusLane[57][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane22_strm0_data_valid    ( DownstreamStackBusLane[57][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane22_strm1_ready         ( DownstreamStackBusLane[57][22].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane22_strm1_cntl          ( DownstreamStackBusLane[57][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane22_strm1_data          ( DownstreamStackBusLane[57][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane22_strm1_data_valid    ( DownstreamStackBusLane[57][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane23_strm0_ready         ( DownstreamStackBusLane[57][23].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane23_strm0_cntl          ( DownstreamStackBusLane[57][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane23_strm0_data          ( DownstreamStackBusLane[57][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane23_strm0_data_valid    ( DownstreamStackBusLane[57][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane23_strm1_ready         ( DownstreamStackBusLane[57][23].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane23_strm1_cntl          ( DownstreamStackBusLane[57][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane23_strm1_data          ( DownstreamStackBusLane[57][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane23_strm1_data_valid    ( DownstreamStackBusLane[57][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane24_strm0_ready         ( DownstreamStackBusLane[57][24].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane24_strm0_cntl          ( DownstreamStackBusLane[57][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane24_strm0_data          ( DownstreamStackBusLane[57][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane24_strm0_data_valid    ( DownstreamStackBusLane[57][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane24_strm1_ready         ( DownstreamStackBusLane[57][24].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane24_strm1_cntl          ( DownstreamStackBusLane[57][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane24_strm1_data          ( DownstreamStackBusLane[57][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane24_strm1_data_valid    ( DownstreamStackBusLane[57][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane25_strm0_ready         ( DownstreamStackBusLane[57][25].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane25_strm0_cntl          ( DownstreamStackBusLane[57][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane25_strm0_data          ( DownstreamStackBusLane[57][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane25_strm0_data_valid    ( DownstreamStackBusLane[57][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane25_strm1_ready         ( DownstreamStackBusLane[57][25].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane25_strm1_cntl          ( DownstreamStackBusLane[57][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane25_strm1_data          ( DownstreamStackBusLane[57][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane25_strm1_data_valid    ( DownstreamStackBusLane[57][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane26_strm0_ready         ( DownstreamStackBusLane[57][26].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane26_strm0_cntl          ( DownstreamStackBusLane[57][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane26_strm0_data          ( DownstreamStackBusLane[57][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane26_strm0_data_valid    ( DownstreamStackBusLane[57][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane26_strm1_ready         ( DownstreamStackBusLane[57][26].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane26_strm1_cntl          ( DownstreamStackBusLane[57][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane26_strm1_data          ( DownstreamStackBusLane[57][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane26_strm1_data_valid    ( DownstreamStackBusLane[57][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane27_strm0_ready         ( DownstreamStackBusLane[57][27].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane27_strm0_cntl          ( DownstreamStackBusLane[57][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane27_strm0_data          ( DownstreamStackBusLane[57][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane27_strm0_data_valid    ( DownstreamStackBusLane[57][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane27_strm1_ready         ( DownstreamStackBusLane[57][27].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane27_strm1_cntl          ( DownstreamStackBusLane[57][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane27_strm1_data          ( DownstreamStackBusLane[57][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane27_strm1_data_valid    ( DownstreamStackBusLane[57][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane28_strm0_ready         ( DownstreamStackBusLane[57][28].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane28_strm0_cntl          ( DownstreamStackBusLane[57][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane28_strm0_data          ( DownstreamStackBusLane[57][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane28_strm0_data_valid    ( DownstreamStackBusLane[57][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane28_strm1_ready         ( DownstreamStackBusLane[57][28].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane28_strm1_cntl          ( DownstreamStackBusLane[57][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane28_strm1_data          ( DownstreamStackBusLane[57][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane28_strm1_data_valid    ( DownstreamStackBusLane[57][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane29_strm0_ready         ( DownstreamStackBusLane[57][29].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane29_strm0_cntl          ( DownstreamStackBusLane[57][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane29_strm0_data          ( DownstreamStackBusLane[57][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane29_strm0_data_valid    ( DownstreamStackBusLane[57][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane29_strm1_ready         ( DownstreamStackBusLane[57][29].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane29_strm1_cntl          ( DownstreamStackBusLane[57][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane29_strm1_data          ( DownstreamStackBusLane[57][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane29_strm1_data_valid    ( DownstreamStackBusLane[57][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane30_strm0_ready         ( DownstreamStackBusLane[57][30].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane30_strm0_cntl          ( DownstreamStackBusLane[57][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane30_strm0_data          ( DownstreamStackBusLane[57][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane30_strm0_data_valid    ( DownstreamStackBusLane[57][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane30_strm1_ready         ( DownstreamStackBusLane[57][30].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane30_strm1_cntl          ( DownstreamStackBusLane[57][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane30_strm1_data          ( DownstreamStackBusLane[57][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane30_strm1_data_valid    ( DownstreamStackBusLane[57][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 57, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane31_strm0_ready         ( DownstreamStackBusLane[57][31].pe__std__lane_strm0_ready              ),      
        .std__pe57__lane31_strm0_cntl          ( DownstreamStackBusLane[57][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe57__lane31_strm0_data          ( DownstreamStackBusLane[57][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe57__lane31_strm0_data_valid    ( DownstreamStackBusLane[57][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__std__lane31_strm1_ready         ( DownstreamStackBusLane[57][31].pe__std__lane_strm1_ready              ),      
        .std__pe57__lane31_strm1_cntl          ( DownstreamStackBusLane[57][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe57__lane31_strm1_data          ( DownstreamStackBusLane[57][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe57__lane31_strm1_data_valid    ( DownstreamStackBusLane[57][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane0_strm0_ready         ( DownstreamStackBusLane[58][0].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane0_strm0_cntl          ( DownstreamStackBusLane[58][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane0_strm0_data          ( DownstreamStackBusLane[58][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane0_strm0_data_valid    ( DownstreamStackBusLane[58][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane0_strm1_ready         ( DownstreamStackBusLane[58][0].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane0_strm1_cntl          ( DownstreamStackBusLane[58][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane0_strm1_data          ( DownstreamStackBusLane[58][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane0_strm1_data_valid    ( DownstreamStackBusLane[58][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane1_strm0_ready         ( DownstreamStackBusLane[58][1].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane1_strm0_cntl          ( DownstreamStackBusLane[58][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane1_strm0_data          ( DownstreamStackBusLane[58][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane1_strm0_data_valid    ( DownstreamStackBusLane[58][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane1_strm1_ready         ( DownstreamStackBusLane[58][1].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane1_strm1_cntl          ( DownstreamStackBusLane[58][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane1_strm1_data          ( DownstreamStackBusLane[58][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane1_strm1_data_valid    ( DownstreamStackBusLane[58][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane2_strm0_ready         ( DownstreamStackBusLane[58][2].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane2_strm0_cntl          ( DownstreamStackBusLane[58][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane2_strm0_data          ( DownstreamStackBusLane[58][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane2_strm0_data_valid    ( DownstreamStackBusLane[58][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane2_strm1_ready         ( DownstreamStackBusLane[58][2].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane2_strm1_cntl          ( DownstreamStackBusLane[58][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane2_strm1_data          ( DownstreamStackBusLane[58][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane2_strm1_data_valid    ( DownstreamStackBusLane[58][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane3_strm0_ready         ( DownstreamStackBusLane[58][3].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane3_strm0_cntl          ( DownstreamStackBusLane[58][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane3_strm0_data          ( DownstreamStackBusLane[58][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane3_strm0_data_valid    ( DownstreamStackBusLane[58][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane3_strm1_ready         ( DownstreamStackBusLane[58][3].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane3_strm1_cntl          ( DownstreamStackBusLane[58][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane3_strm1_data          ( DownstreamStackBusLane[58][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane3_strm1_data_valid    ( DownstreamStackBusLane[58][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane4_strm0_ready         ( DownstreamStackBusLane[58][4].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane4_strm0_cntl          ( DownstreamStackBusLane[58][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane4_strm0_data          ( DownstreamStackBusLane[58][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane4_strm0_data_valid    ( DownstreamStackBusLane[58][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane4_strm1_ready         ( DownstreamStackBusLane[58][4].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane4_strm1_cntl          ( DownstreamStackBusLane[58][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane4_strm1_data          ( DownstreamStackBusLane[58][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane4_strm1_data_valid    ( DownstreamStackBusLane[58][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane5_strm0_ready         ( DownstreamStackBusLane[58][5].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane5_strm0_cntl          ( DownstreamStackBusLane[58][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane5_strm0_data          ( DownstreamStackBusLane[58][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane5_strm0_data_valid    ( DownstreamStackBusLane[58][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane5_strm1_ready         ( DownstreamStackBusLane[58][5].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane5_strm1_cntl          ( DownstreamStackBusLane[58][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane5_strm1_data          ( DownstreamStackBusLane[58][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane5_strm1_data_valid    ( DownstreamStackBusLane[58][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane6_strm0_ready         ( DownstreamStackBusLane[58][6].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane6_strm0_cntl          ( DownstreamStackBusLane[58][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane6_strm0_data          ( DownstreamStackBusLane[58][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane6_strm0_data_valid    ( DownstreamStackBusLane[58][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane6_strm1_ready         ( DownstreamStackBusLane[58][6].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane6_strm1_cntl          ( DownstreamStackBusLane[58][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane6_strm1_data          ( DownstreamStackBusLane[58][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane6_strm1_data_valid    ( DownstreamStackBusLane[58][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane7_strm0_ready         ( DownstreamStackBusLane[58][7].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane7_strm0_cntl          ( DownstreamStackBusLane[58][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane7_strm0_data          ( DownstreamStackBusLane[58][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane7_strm0_data_valid    ( DownstreamStackBusLane[58][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane7_strm1_ready         ( DownstreamStackBusLane[58][7].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane7_strm1_cntl          ( DownstreamStackBusLane[58][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane7_strm1_data          ( DownstreamStackBusLane[58][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane7_strm1_data_valid    ( DownstreamStackBusLane[58][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane8_strm0_ready         ( DownstreamStackBusLane[58][8].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane8_strm0_cntl          ( DownstreamStackBusLane[58][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane8_strm0_data          ( DownstreamStackBusLane[58][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane8_strm0_data_valid    ( DownstreamStackBusLane[58][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane8_strm1_ready         ( DownstreamStackBusLane[58][8].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane8_strm1_cntl          ( DownstreamStackBusLane[58][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane8_strm1_data          ( DownstreamStackBusLane[58][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane8_strm1_data_valid    ( DownstreamStackBusLane[58][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane9_strm0_ready         ( DownstreamStackBusLane[58][9].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane9_strm0_cntl          ( DownstreamStackBusLane[58][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane9_strm0_data          ( DownstreamStackBusLane[58][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane9_strm0_data_valid    ( DownstreamStackBusLane[58][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane9_strm1_ready         ( DownstreamStackBusLane[58][9].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane9_strm1_cntl          ( DownstreamStackBusLane[58][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane9_strm1_data          ( DownstreamStackBusLane[58][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane9_strm1_data_valid    ( DownstreamStackBusLane[58][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane10_strm0_ready         ( DownstreamStackBusLane[58][10].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane10_strm0_cntl          ( DownstreamStackBusLane[58][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane10_strm0_data          ( DownstreamStackBusLane[58][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane10_strm0_data_valid    ( DownstreamStackBusLane[58][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane10_strm1_ready         ( DownstreamStackBusLane[58][10].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane10_strm1_cntl          ( DownstreamStackBusLane[58][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane10_strm1_data          ( DownstreamStackBusLane[58][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane10_strm1_data_valid    ( DownstreamStackBusLane[58][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane11_strm0_ready         ( DownstreamStackBusLane[58][11].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane11_strm0_cntl          ( DownstreamStackBusLane[58][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane11_strm0_data          ( DownstreamStackBusLane[58][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane11_strm0_data_valid    ( DownstreamStackBusLane[58][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane11_strm1_ready         ( DownstreamStackBusLane[58][11].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane11_strm1_cntl          ( DownstreamStackBusLane[58][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane11_strm1_data          ( DownstreamStackBusLane[58][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane11_strm1_data_valid    ( DownstreamStackBusLane[58][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane12_strm0_ready         ( DownstreamStackBusLane[58][12].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane12_strm0_cntl          ( DownstreamStackBusLane[58][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane12_strm0_data          ( DownstreamStackBusLane[58][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane12_strm0_data_valid    ( DownstreamStackBusLane[58][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane12_strm1_ready         ( DownstreamStackBusLane[58][12].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane12_strm1_cntl          ( DownstreamStackBusLane[58][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane12_strm1_data          ( DownstreamStackBusLane[58][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane12_strm1_data_valid    ( DownstreamStackBusLane[58][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane13_strm0_ready         ( DownstreamStackBusLane[58][13].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane13_strm0_cntl          ( DownstreamStackBusLane[58][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane13_strm0_data          ( DownstreamStackBusLane[58][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane13_strm0_data_valid    ( DownstreamStackBusLane[58][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane13_strm1_ready         ( DownstreamStackBusLane[58][13].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane13_strm1_cntl          ( DownstreamStackBusLane[58][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane13_strm1_data          ( DownstreamStackBusLane[58][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane13_strm1_data_valid    ( DownstreamStackBusLane[58][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane14_strm0_ready         ( DownstreamStackBusLane[58][14].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane14_strm0_cntl          ( DownstreamStackBusLane[58][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane14_strm0_data          ( DownstreamStackBusLane[58][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane14_strm0_data_valid    ( DownstreamStackBusLane[58][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane14_strm1_ready         ( DownstreamStackBusLane[58][14].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane14_strm1_cntl          ( DownstreamStackBusLane[58][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane14_strm1_data          ( DownstreamStackBusLane[58][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane14_strm1_data_valid    ( DownstreamStackBusLane[58][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane15_strm0_ready         ( DownstreamStackBusLane[58][15].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane15_strm0_cntl          ( DownstreamStackBusLane[58][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane15_strm0_data          ( DownstreamStackBusLane[58][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane15_strm0_data_valid    ( DownstreamStackBusLane[58][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane15_strm1_ready         ( DownstreamStackBusLane[58][15].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane15_strm1_cntl          ( DownstreamStackBusLane[58][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane15_strm1_data          ( DownstreamStackBusLane[58][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane15_strm1_data_valid    ( DownstreamStackBusLane[58][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane16_strm0_ready         ( DownstreamStackBusLane[58][16].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane16_strm0_cntl          ( DownstreamStackBusLane[58][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane16_strm0_data          ( DownstreamStackBusLane[58][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane16_strm0_data_valid    ( DownstreamStackBusLane[58][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane16_strm1_ready         ( DownstreamStackBusLane[58][16].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane16_strm1_cntl          ( DownstreamStackBusLane[58][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane16_strm1_data          ( DownstreamStackBusLane[58][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane16_strm1_data_valid    ( DownstreamStackBusLane[58][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane17_strm0_ready         ( DownstreamStackBusLane[58][17].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane17_strm0_cntl          ( DownstreamStackBusLane[58][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane17_strm0_data          ( DownstreamStackBusLane[58][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane17_strm0_data_valid    ( DownstreamStackBusLane[58][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane17_strm1_ready         ( DownstreamStackBusLane[58][17].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane17_strm1_cntl          ( DownstreamStackBusLane[58][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane17_strm1_data          ( DownstreamStackBusLane[58][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane17_strm1_data_valid    ( DownstreamStackBusLane[58][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane18_strm0_ready         ( DownstreamStackBusLane[58][18].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane18_strm0_cntl          ( DownstreamStackBusLane[58][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane18_strm0_data          ( DownstreamStackBusLane[58][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane18_strm0_data_valid    ( DownstreamStackBusLane[58][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane18_strm1_ready         ( DownstreamStackBusLane[58][18].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane18_strm1_cntl          ( DownstreamStackBusLane[58][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane18_strm1_data          ( DownstreamStackBusLane[58][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane18_strm1_data_valid    ( DownstreamStackBusLane[58][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane19_strm0_ready         ( DownstreamStackBusLane[58][19].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane19_strm0_cntl          ( DownstreamStackBusLane[58][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane19_strm0_data          ( DownstreamStackBusLane[58][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane19_strm0_data_valid    ( DownstreamStackBusLane[58][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane19_strm1_ready         ( DownstreamStackBusLane[58][19].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane19_strm1_cntl          ( DownstreamStackBusLane[58][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane19_strm1_data          ( DownstreamStackBusLane[58][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane19_strm1_data_valid    ( DownstreamStackBusLane[58][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane20_strm0_ready         ( DownstreamStackBusLane[58][20].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane20_strm0_cntl          ( DownstreamStackBusLane[58][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane20_strm0_data          ( DownstreamStackBusLane[58][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane20_strm0_data_valid    ( DownstreamStackBusLane[58][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane20_strm1_ready         ( DownstreamStackBusLane[58][20].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane20_strm1_cntl          ( DownstreamStackBusLane[58][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane20_strm1_data          ( DownstreamStackBusLane[58][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane20_strm1_data_valid    ( DownstreamStackBusLane[58][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane21_strm0_ready         ( DownstreamStackBusLane[58][21].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane21_strm0_cntl          ( DownstreamStackBusLane[58][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane21_strm0_data          ( DownstreamStackBusLane[58][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane21_strm0_data_valid    ( DownstreamStackBusLane[58][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane21_strm1_ready         ( DownstreamStackBusLane[58][21].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane21_strm1_cntl          ( DownstreamStackBusLane[58][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane21_strm1_data          ( DownstreamStackBusLane[58][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane21_strm1_data_valid    ( DownstreamStackBusLane[58][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane22_strm0_ready         ( DownstreamStackBusLane[58][22].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane22_strm0_cntl          ( DownstreamStackBusLane[58][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane22_strm0_data          ( DownstreamStackBusLane[58][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane22_strm0_data_valid    ( DownstreamStackBusLane[58][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane22_strm1_ready         ( DownstreamStackBusLane[58][22].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane22_strm1_cntl          ( DownstreamStackBusLane[58][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane22_strm1_data          ( DownstreamStackBusLane[58][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane22_strm1_data_valid    ( DownstreamStackBusLane[58][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane23_strm0_ready         ( DownstreamStackBusLane[58][23].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane23_strm0_cntl          ( DownstreamStackBusLane[58][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane23_strm0_data          ( DownstreamStackBusLane[58][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane23_strm0_data_valid    ( DownstreamStackBusLane[58][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane23_strm1_ready         ( DownstreamStackBusLane[58][23].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane23_strm1_cntl          ( DownstreamStackBusLane[58][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane23_strm1_data          ( DownstreamStackBusLane[58][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane23_strm1_data_valid    ( DownstreamStackBusLane[58][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane24_strm0_ready         ( DownstreamStackBusLane[58][24].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane24_strm0_cntl          ( DownstreamStackBusLane[58][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane24_strm0_data          ( DownstreamStackBusLane[58][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane24_strm0_data_valid    ( DownstreamStackBusLane[58][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane24_strm1_ready         ( DownstreamStackBusLane[58][24].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane24_strm1_cntl          ( DownstreamStackBusLane[58][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane24_strm1_data          ( DownstreamStackBusLane[58][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane24_strm1_data_valid    ( DownstreamStackBusLane[58][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane25_strm0_ready         ( DownstreamStackBusLane[58][25].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane25_strm0_cntl          ( DownstreamStackBusLane[58][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane25_strm0_data          ( DownstreamStackBusLane[58][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane25_strm0_data_valid    ( DownstreamStackBusLane[58][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane25_strm1_ready         ( DownstreamStackBusLane[58][25].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane25_strm1_cntl          ( DownstreamStackBusLane[58][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane25_strm1_data          ( DownstreamStackBusLane[58][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane25_strm1_data_valid    ( DownstreamStackBusLane[58][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane26_strm0_ready         ( DownstreamStackBusLane[58][26].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane26_strm0_cntl          ( DownstreamStackBusLane[58][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane26_strm0_data          ( DownstreamStackBusLane[58][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane26_strm0_data_valid    ( DownstreamStackBusLane[58][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane26_strm1_ready         ( DownstreamStackBusLane[58][26].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane26_strm1_cntl          ( DownstreamStackBusLane[58][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane26_strm1_data          ( DownstreamStackBusLane[58][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane26_strm1_data_valid    ( DownstreamStackBusLane[58][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane27_strm0_ready         ( DownstreamStackBusLane[58][27].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane27_strm0_cntl          ( DownstreamStackBusLane[58][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane27_strm0_data          ( DownstreamStackBusLane[58][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane27_strm0_data_valid    ( DownstreamStackBusLane[58][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane27_strm1_ready         ( DownstreamStackBusLane[58][27].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane27_strm1_cntl          ( DownstreamStackBusLane[58][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane27_strm1_data          ( DownstreamStackBusLane[58][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane27_strm1_data_valid    ( DownstreamStackBusLane[58][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane28_strm0_ready         ( DownstreamStackBusLane[58][28].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane28_strm0_cntl          ( DownstreamStackBusLane[58][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane28_strm0_data          ( DownstreamStackBusLane[58][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane28_strm0_data_valid    ( DownstreamStackBusLane[58][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane28_strm1_ready         ( DownstreamStackBusLane[58][28].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane28_strm1_cntl          ( DownstreamStackBusLane[58][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane28_strm1_data          ( DownstreamStackBusLane[58][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane28_strm1_data_valid    ( DownstreamStackBusLane[58][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane29_strm0_ready         ( DownstreamStackBusLane[58][29].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane29_strm0_cntl          ( DownstreamStackBusLane[58][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane29_strm0_data          ( DownstreamStackBusLane[58][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane29_strm0_data_valid    ( DownstreamStackBusLane[58][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane29_strm1_ready         ( DownstreamStackBusLane[58][29].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane29_strm1_cntl          ( DownstreamStackBusLane[58][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane29_strm1_data          ( DownstreamStackBusLane[58][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane29_strm1_data_valid    ( DownstreamStackBusLane[58][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane30_strm0_ready         ( DownstreamStackBusLane[58][30].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane30_strm0_cntl          ( DownstreamStackBusLane[58][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane30_strm0_data          ( DownstreamStackBusLane[58][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane30_strm0_data_valid    ( DownstreamStackBusLane[58][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane30_strm1_ready         ( DownstreamStackBusLane[58][30].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane30_strm1_cntl          ( DownstreamStackBusLane[58][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane30_strm1_data          ( DownstreamStackBusLane[58][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane30_strm1_data_valid    ( DownstreamStackBusLane[58][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 58, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane31_strm0_ready         ( DownstreamStackBusLane[58][31].pe__std__lane_strm0_ready              ),      
        .std__pe58__lane31_strm0_cntl          ( DownstreamStackBusLane[58][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe58__lane31_strm0_data          ( DownstreamStackBusLane[58][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe58__lane31_strm0_data_valid    ( DownstreamStackBusLane[58][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__std__lane31_strm1_ready         ( DownstreamStackBusLane[58][31].pe__std__lane_strm1_ready              ),      
        .std__pe58__lane31_strm1_cntl          ( DownstreamStackBusLane[58][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe58__lane31_strm1_data          ( DownstreamStackBusLane[58][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe58__lane31_strm1_data_valid    ( DownstreamStackBusLane[58][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane0_strm0_ready         ( DownstreamStackBusLane[59][0].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane0_strm0_cntl          ( DownstreamStackBusLane[59][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane0_strm0_data          ( DownstreamStackBusLane[59][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane0_strm0_data_valid    ( DownstreamStackBusLane[59][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane0_strm1_ready         ( DownstreamStackBusLane[59][0].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane0_strm1_cntl          ( DownstreamStackBusLane[59][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane0_strm1_data          ( DownstreamStackBusLane[59][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane0_strm1_data_valid    ( DownstreamStackBusLane[59][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane1_strm0_ready         ( DownstreamStackBusLane[59][1].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane1_strm0_cntl          ( DownstreamStackBusLane[59][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane1_strm0_data          ( DownstreamStackBusLane[59][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane1_strm0_data_valid    ( DownstreamStackBusLane[59][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane1_strm1_ready         ( DownstreamStackBusLane[59][1].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane1_strm1_cntl          ( DownstreamStackBusLane[59][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane1_strm1_data          ( DownstreamStackBusLane[59][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane1_strm1_data_valid    ( DownstreamStackBusLane[59][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane2_strm0_ready         ( DownstreamStackBusLane[59][2].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane2_strm0_cntl          ( DownstreamStackBusLane[59][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane2_strm0_data          ( DownstreamStackBusLane[59][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane2_strm0_data_valid    ( DownstreamStackBusLane[59][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane2_strm1_ready         ( DownstreamStackBusLane[59][2].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane2_strm1_cntl          ( DownstreamStackBusLane[59][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane2_strm1_data          ( DownstreamStackBusLane[59][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane2_strm1_data_valid    ( DownstreamStackBusLane[59][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane3_strm0_ready         ( DownstreamStackBusLane[59][3].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane3_strm0_cntl          ( DownstreamStackBusLane[59][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane3_strm0_data          ( DownstreamStackBusLane[59][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane3_strm0_data_valid    ( DownstreamStackBusLane[59][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane3_strm1_ready         ( DownstreamStackBusLane[59][3].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane3_strm1_cntl          ( DownstreamStackBusLane[59][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane3_strm1_data          ( DownstreamStackBusLane[59][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane3_strm1_data_valid    ( DownstreamStackBusLane[59][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane4_strm0_ready         ( DownstreamStackBusLane[59][4].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane4_strm0_cntl          ( DownstreamStackBusLane[59][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane4_strm0_data          ( DownstreamStackBusLane[59][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane4_strm0_data_valid    ( DownstreamStackBusLane[59][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane4_strm1_ready         ( DownstreamStackBusLane[59][4].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane4_strm1_cntl          ( DownstreamStackBusLane[59][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane4_strm1_data          ( DownstreamStackBusLane[59][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane4_strm1_data_valid    ( DownstreamStackBusLane[59][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane5_strm0_ready         ( DownstreamStackBusLane[59][5].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane5_strm0_cntl          ( DownstreamStackBusLane[59][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane5_strm0_data          ( DownstreamStackBusLane[59][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane5_strm0_data_valid    ( DownstreamStackBusLane[59][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane5_strm1_ready         ( DownstreamStackBusLane[59][5].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane5_strm1_cntl          ( DownstreamStackBusLane[59][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane5_strm1_data          ( DownstreamStackBusLane[59][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane5_strm1_data_valid    ( DownstreamStackBusLane[59][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane6_strm0_ready         ( DownstreamStackBusLane[59][6].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane6_strm0_cntl          ( DownstreamStackBusLane[59][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane6_strm0_data          ( DownstreamStackBusLane[59][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane6_strm0_data_valid    ( DownstreamStackBusLane[59][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane6_strm1_ready         ( DownstreamStackBusLane[59][6].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane6_strm1_cntl          ( DownstreamStackBusLane[59][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane6_strm1_data          ( DownstreamStackBusLane[59][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane6_strm1_data_valid    ( DownstreamStackBusLane[59][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane7_strm0_ready         ( DownstreamStackBusLane[59][7].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane7_strm0_cntl          ( DownstreamStackBusLane[59][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane7_strm0_data          ( DownstreamStackBusLane[59][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane7_strm0_data_valid    ( DownstreamStackBusLane[59][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane7_strm1_ready         ( DownstreamStackBusLane[59][7].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane7_strm1_cntl          ( DownstreamStackBusLane[59][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane7_strm1_data          ( DownstreamStackBusLane[59][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane7_strm1_data_valid    ( DownstreamStackBusLane[59][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane8_strm0_ready         ( DownstreamStackBusLane[59][8].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane8_strm0_cntl          ( DownstreamStackBusLane[59][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane8_strm0_data          ( DownstreamStackBusLane[59][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane8_strm0_data_valid    ( DownstreamStackBusLane[59][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane8_strm1_ready         ( DownstreamStackBusLane[59][8].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane8_strm1_cntl          ( DownstreamStackBusLane[59][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane8_strm1_data          ( DownstreamStackBusLane[59][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane8_strm1_data_valid    ( DownstreamStackBusLane[59][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane9_strm0_ready         ( DownstreamStackBusLane[59][9].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane9_strm0_cntl          ( DownstreamStackBusLane[59][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane9_strm0_data          ( DownstreamStackBusLane[59][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane9_strm0_data_valid    ( DownstreamStackBusLane[59][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane9_strm1_ready         ( DownstreamStackBusLane[59][9].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane9_strm1_cntl          ( DownstreamStackBusLane[59][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane9_strm1_data          ( DownstreamStackBusLane[59][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane9_strm1_data_valid    ( DownstreamStackBusLane[59][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane10_strm0_ready         ( DownstreamStackBusLane[59][10].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane10_strm0_cntl          ( DownstreamStackBusLane[59][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane10_strm0_data          ( DownstreamStackBusLane[59][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane10_strm0_data_valid    ( DownstreamStackBusLane[59][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane10_strm1_ready         ( DownstreamStackBusLane[59][10].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane10_strm1_cntl          ( DownstreamStackBusLane[59][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane10_strm1_data          ( DownstreamStackBusLane[59][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane10_strm1_data_valid    ( DownstreamStackBusLane[59][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane11_strm0_ready         ( DownstreamStackBusLane[59][11].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane11_strm0_cntl          ( DownstreamStackBusLane[59][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane11_strm0_data          ( DownstreamStackBusLane[59][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane11_strm0_data_valid    ( DownstreamStackBusLane[59][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane11_strm1_ready         ( DownstreamStackBusLane[59][11].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane11_strm1_cntl          ( DownstreamStackBusLane[59][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane11_strm1_data          ( DownstreamStackBusLane[59][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane11_strm1_data_valid    ( DownstreamStackBusLane[59][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane12_strm0_ready         ( DownstreamStackBusLane[59][12].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane12_strm0_cntl          ( DownstreamStackBusLane[59][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane12_strm0_data          ( DownstreamStackBusLane[59][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane12_strm0_data_valid    ( DownstreamStackBusLane[59][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane12_strm1_ready         ( DownstreamStackBusLane[59][12].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane12_strm1_cntl          ( DownstreamStackBusLane[59][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane12_strm1_data          ( DownstreamStackBusLane[59][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane12_strm1_data_valid    ( DownstreamStackBusLane[59][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane13_strm0_ready         ( DownstreamStackBusLane[59][13].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane13_strm0_cntl          ( DownstreamStackBusLane[59][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane13_strm0_data          ( DownstreamStackBusLane[59][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane13_strm0_data_valid    ( DownstreamStackBusLane[59][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane13_strm1_ready         ( DownstreamStackBusLane[59][13].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane13_strm1_cntl          ( DownstreamStackBusLane[59][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane13_strm1_data          ( DownstreamStackBusLane[59][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane13_strm1_data_valid    ( DownstreamStackBusLane[59][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane14_strm0_ready         ( DownstreamStackBusLane[59][14].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane14_strm0_cntl          ( DownstreamStackBusLane[59][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane14_strm0_data          ( DownstreamStackBusLane[59][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane14_strm0_data_valid    ( DownstreamStackBusLane[59][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane14_strm1_ready         ( DownstreamStackBusLane[59][14].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane14_strm1_cntl          ( DownstreamStackBusLane[59][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane14_strm1_data          ( DownstreamStackBusLane[59][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane14_strm1_data_valid    ( DownstreamStackBusLane[59][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane15_strm0_ready         ( DownstreamStackBusLane[59][15].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane15_strm0_cntl          ( DownstreamStackBusLane[59][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane15_strm0_data          ( DownstreamStackBusLane[59][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane15_strm0_data_valid    ( DownstreamStackBusLane[59][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane15_strm1_ready         ( DownstreamStackBusLane[59][15].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane15_strm1_cntl          ( DownstreamStackBusLane[59][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane15_strm1_data          ( DownstreamStackBusLane[59][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane15_strm1_data_valid    ( DownstreamStackBusLane[59][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane16_strm0_ready         ( DownstreamStackBusLane[59][16].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane16_strm0_cntl          ( DownstreamStackBusLane[59][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane16_strm0_data          ( DownstreamStackBusLane[59][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane16_strm0_data_valid    ( DownstreamStackBusLane[59][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane16_strm1_ready         ( DownstreamStackBusLane[59][16].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane16_strm1_cntl          ( DownstreamStackBusLane[59][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane16_strm1_data          ( DownstreamStackBusLane[59][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane16_strm1_data_valid    ( DownstreamStackBusLane[59][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane17_strm0_ready         ( DownstreamStackBusLane[59][17].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane17_strm0_cntl          ( DownstreamStackBusLane[59][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane17_strm0_data          ( DownstreamStackBusLane[59][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane17_strm0_data_valid    ( DownstreamStackBusLane[59][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane17_strm1_ready         ( DownstreamStackBusLane[59][17].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane17_strm1_cntl          ( DownstreamStackBusLane[59][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane17_strm1_data          ( DownstreamStackBusLane[59][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane17_strm1_data_valid    ( DownstreamStackBusLane[59][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane18_strm0_ready         ( DownstreamStackBusLane[59][18].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane18_strm0_cntl          ( DownstreamStackBusLane[59][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane18_strm0_data          ( DownstreamStackBusLane[59][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane18_strm0_data_valid    ( DownstreamStackBusLane[59][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane18_strm1_ready         ( DownstreamStackBusLane[59][18].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane18_strm1_cntl          ( DownstreamStackBusLane[59][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane18_strm1_data          ( DownstreamStackBusLane[59][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane18_strm1_data_valid    ( DownstreamStackBusLane[59][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane19_strm0_ready         ( DownstreamStackBusLane[59][19].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane19_strm0_cntl          ( DownstreamStackBusLane[59][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane19_strm0_data          ( DownstreamStackBusLane[59][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane19_strm0_data_valid    ( DownstreamStackBusLane[59][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane19_strm1_ready         ( DownstreamStackBusLane[59][19].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane19_strm1_cntl          ( DownstreamStackBusLane[59][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane19_strm1_data          ( DownstreamStackBusLane[59][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane19_strm1_data_valid    ( DownstreamStackBusLane[59][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane20_strm0_ready         ( DownstreamStackBusLane[59][20].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane20_strm0_cntl          ( DownstreamStackBusLane[59][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane20_strm0_data          ( DownstreamStackBusLane[59][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane20_strm0_data_valid    ( DownstreamStackBusLane[59][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane20_strm1_ready         ( DownstreamStackBusLane[59][20].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane20_strm1_cntl          ( DownstreamStackBusLane[59][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane20_strm1_data          ( DownstreamStackBusLane[59][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane20_strm1_data_valid    ( DownstreamStackBusLane[59][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane21_strm0_ready         ( DownstreamStackBusLane[59][21].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane21_strm0_cntl          ( DownstreamStackBusLane[59][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane21_strm0_data          ( DownstreamStackBusLane[59][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane21_strm0_data_valid    ( DownstreamStackBusLane[59][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane21_strm1_ready         ( DownstreamStackBusLane[59][21].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane21_strm1_cntl          ( DownstreamStackBusLane[59][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane21_strm1_data          ( DownstreamStackBusLane[59][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane21_strm1_data_valid    ( DownstreamStackBusLane[59][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane22_strm0_ready         ( DownstreamStackBusLane[59][22].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane22_strm0_cntl          ( DownstreamStackBusLane[59][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane22_strm0_data          ( DownstreamStackBusLane[59][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane22_strm0_data_valid    ( DownstreamStackBusLane[59][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane22_strm1_ready         ( DownstreamStackBusLane[59][22].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane22_strm1_cntl          ( DownstreamStackBusLane[59][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane22_strm1_data          ( DownstreamStackBusLane[59][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane22_strm1_data_valid    ( DownstreamStackBusLane[59][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane23_strm0_ready         ( DownstreamStackBusLane[59][23].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane23_strm0_cntl          ( DownstreamStackBusLane[59][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane23_strm0_data          ( DownstreamStackBusLane[59][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane23_strm0_data_valid    ( DownstreamStackBusLane[59][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane23_strm1_ready         ( DownstreamStackBusLane[59][23].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane23_strm1_cntl          ( DownstreamStackBusLane[59][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane23_strm1_data          ( DownstreamStackBusLane[59][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane23_strm1_data_valid    ( DownstreamStackBusLane[59][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane24_strm0_ready         ( DownstreamStackBusLane[59][24].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane24_strm0_cntl          ( DownstreamStackBusLane[59][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane24_strm0_data          ( DownstreamStackBusLane[59][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane24_strm0_data_valid    ( DownstreamStackBusLane[59][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane24_strm1_ready         ( DownstreamStackBusLane[59][24].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane24_strm1_cntl          ( DownstreamStackBusLane[59][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane24_strm1_data          ( DownstreamStackBusLane[59][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane24_strm1_data_valid    ( DownstreamStackBusLane[59][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane25_strm0_ready         ( DownstreamStackBusLane[59][25].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane25_strm0_cntl          ( DownstreamStackBusLane[59][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane25_strm0_data          ( DownstreamStackBusLane[59][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane25_strm0_data_valid    ( DownstreamStackBusLane[59][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane25_strm1_ready         ( DownstreamStackBusLane[59][25].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane25_strm1_cntl          ( DownstreamStackBusLane[59][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane25_strm1_data          ( DownstreamStackBusLane[59][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane25_strm1_data_valid    ( DownstreamStackBusLane[59][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane26_strm0_ready         ( DownstreamStackBusLane[59][26].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane26_strm0_cntl          ( DownstreamStackBusLane[59][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane26_strm0_data          ( DownstreamStackBusLane[59][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane26_strm0_data_valid    ( DownstreamStackBusLane[59][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane26_strm1_ready         ( DownstreamStackBusLane[59][26].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane26_strm1_cntl          ( DownstreamStackBusLane[59][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane26_strm1_data          ( DownstreamStackBusLane[59][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane26_strm1_data_valid    ( DownstreamStackBusLane[59][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane27_strm0_ready         ( DownstreamStackBusLane[59][27].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane27_strm0_cntl          ( DownstreamStackBusLane[59][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane27_strm0_data          ( DownstreamStackBusLane[59][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane27_strm0_data_valid    ( DownstreamStackBusLane[59][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane27_strm1_ready         ( DownstreamStackBusLane[59][27].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane27_strm1_cntl          ( DownstreamStackBusLane[59][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane27_strm1_data          ( DownstreamStackBusLane[59][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane27_strm1_data_valid    ( DownstreamStackBusLane[59][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane28_strm0_ready         ( DownstreamStackBusLane[59][28].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane28_strm0_cntl          ( DownstreamStackBusLane[59][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane28_strm0_data          ( DownstreamStackBusLane[59][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane28_strm0_data_valid    ( DownstreamStackBusLane[59][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane28_strm1_ready         ( DownstreamStackBusLane[59][28].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane28_strm1_cntl          ( DownstreamStackBusLane[59][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane28_strm1_data          ( DownstreamStackBusLane[59][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane28_strm1_data_valid    ( DownstreamStackBusLane[59][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane29_strm0_ready         ( DownstreamStackBusLane[59][29].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane29_strm0_cntl          ( DownstreamStackBusLane[59][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane29_strm0_data          ( DownstreamStackBusLane[59][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane29_strm0_data_valid    ( DownstreamStackBusLane[59][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane29_strm1_ready         ( DownstreamStackBusLane[59][29].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane29_strm1_cntl          ( DownstreamStackBusLane[59][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane29_strm1_data          ( DownstreamStackBusLane[59][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane29_strm1_data_valid    ( DownstreamStackBusLane[59][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane30_strm0_ready         ( DownstreamStackBusLane[59][30].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane30_strm0_cntl          ( DownstreamStackBusLane[59][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane30_strm0_data          ( DownstreamStackBusLane[59][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane30_strm0_data_valid    ( DownstreamStackBusLane[59][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane30_strm1_ready         ( DownstreamStackBusLane[59][30].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane30_strm1_cntl          ( DownstreamStackBusLane[59][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane30_strm1_data          ( DownstreamStackBusLane[59][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane30_strm1_data_valid    ( DownstreamStackBusLane[59][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 59, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane31_strm0_ready         ( DownstreamStackBusLane[59][31].pe__std__lane_strm0_ready              ),      
        .std__pe59__lane31_strm0_cntl          ( DownstreamStackBusLane[59][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe59__lane31_strm0_data          ( DownstreamStackBusLane[59][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe59__lane31_strm0_data_valid    ( DownstreamStackBusLane[59][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__std__lane31_strm1_ready         ( DownstreamStackBusLane[59][31].pe__std__lane_strm1_ready              ),      
        .std__pe59__lane31_strm1_cntl          ( DownstreamStackBusLane[59][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe59__lane31_strm1_data          ( DownstreamStackBusLane[59][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe59__lane31_strm1_data_valid    ( DownstreamStackBusLane[59][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane0_strm0_ready         ( DownstreamStackBusLane[60][0].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane0_strm0_cntl          ( DownstreamStackBusLane[60][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane0_strm0_data          ( DownstreamStackBusLane[60][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane0_strm0_data_valid    ( DownstreamStackBusLane[60][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane0_strm1_ready         ( DownstreamStackBusLane[60][0].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane0_strm1_cntl          ( DownstreamStackBusLane[60][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane0_strm1_data          ( DownstreamStackBusLane[60][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane0_strm1_data_valid    ( DownstreamStackBusLane[60][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane1_strm0_ready         ( DownstreamStackBusLane[60][1].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane1_strm0_cntl          ( DownstreamStackBusLane[60][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane1_strm0_data          ( DownstreamStackBusLane[60][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane1_strm0_data_valid    ( DownstreamStackBusLane[60][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane1_strm1_ready         ( DownstreamStackBusLane[60][1].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane1_strm1_cntl          ( DownstreamStackBusLane[60][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane1_strm1_data          ( DownstreamStackBusLane[60][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane1_strm1_data_valid    ( DownstreamStackBusLane[60][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane2_strm0_ready         ( DownstreamStackBusLane[60][2].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane2_strm0_cntl          ( DownstreamStackBusLane[60][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane2_strm0_data          ( DownstreamStackBusLane[60][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane2_strm0_data_valid    ( DownstreamStackBusLane[60][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane2_strm1_ready         ( DownstreamStackBusLane[60][2].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane2_strm1_cntl          ( DownstreamStackBusLane[60][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane2_strm1_data          ( DownstreamStackBusLane[60][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane2_strm1_data_valid    ( DownstreamStackBusLane[60][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane3_strm0_ready         ( DownstreamStackBusLane[60][3].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane3_strm0_cntl          ( DownstreamStackBusLane[60][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane3_strm0_data          ( DownstreamStackBusLane[60][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane3_strm0_data_valid    ( DownstreamStackBusLane[60][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane3_strm1_ready         ( DownstreamStackBusLane[60][3].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane3_strm1_cntl          ( DownstreamStackBusLane[60][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane3_strm1_data          ( DownstreamStackBusLane[60][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane3_strm1_data_valid    ( DownstreamStackBusLane[60][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane4_strm0_ready         ( DownstreamStackBusLane[60][4].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane4_strm0_cntl          ( DownstreamStackBusLane[60][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane4_strm0_data          ( DownstreamStackBusLane[60][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane4_strm0_data_valid    ( DownstreamStackBusLane[60][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane4_strm1_ready         ( DownstreamStackBusLane[60][4].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane4_strm1_cntl          ( DownstreamStackBusLane[60][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane4_strm1_data          ( DownstreamStackBusLane[60][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane4_strm1_data_valid    ( DownstreamStackBusLane[60][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane5_strm0_ready         ( DownstreamStackBusLane[60][5].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane5_strm0_cntl          ( DownstreamStackBusLane[60][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane5_strm0_data          ( DownstreamStackBusLane[60][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane5_strm0_data_valid    ( DownstreamStackBusLane[60][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane5_strm1_ready         ( DownstreamStackBusLane[60][5].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane5_strm1_cntl          ( DownstreamStackBusLane[60][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane5_strm1_data          ( DownstreamStackBusLane[60][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane5_strm1_data_valid    ( DownstreamStackBusLane[60][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane6_strm0_ready         ( DownstreamStackBusLane[60][6].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane6_strm0_cntl          ( DownstreamStackBusLane[60][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane6_strm0_data          ( DownstreamStackBusLane[60][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane6_strm0_data_valid    ( DownstreamStackBusLane[60][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane6_strm1_ready         ( DownstreamStackBusLane[60][6].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane6_strm1_cntl          ( DownstreamStackBusLane[60][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane6_strm1_data          ( DownstreamStackBusLane[60][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane6_strm1_data_valid    ( DownstreamStackBusLane[60][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane7_strm0_ready         ( DownstreamStackBusLane[60][7].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane7_strm0_cntl          ( DownstreamStackBusLane[60][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane7_strm0_data          ( DownstreamStackBusLane[60][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane7_strm0_data_valid    ( DownstreamStackBusLane[60][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane7_strm1_ready         ( DownstreamStackBusLane[60][7].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane7_strm1_cntl          ( DownstreamStackBusLane[60][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane7_strm1_data          ( DownstreamStackBusLane[60][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane7_strm1_data_valid    ( DownstreamStackBusLane[60][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane8_strm0_ready         ( DownstreamStackBusLane[60][8].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane8_strm0_cntl          ( DownstreamStackBusLane[60][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane8_strm0_data          ( DownstreamStackBusLane[60][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane8_strm0_data_valid    ( DownstreamStackBusLane[60][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane8_strm1_ready         ( DownstreamStackBusLane[60][8].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane8_strm1_cntl          ( DownstreamStackBusLane[60][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane8_strm1_data          ( DownstreamStackBusLane[60][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane8_strm1_data_valid    ( DownstreamStackBusLane[60][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane9_strm0_ready         ( DownstreamStackBusLane[60][9].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane9_strm0_cntl          ( DownstreamStackBusLane[60][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane9_strm0_data          ( DownstreamStackBusLane[60][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane9_strm0_data_valid    ( DownstreamStackBusLane[60][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane9_strm1_ready         ( DownstreamStackBusLane[60][9].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane9_strm1_cntl          ( DownstreamStackBusLane[60][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane9_strm1_data          ( DownstreamStackBusLane[60][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane9_strm1_data_valid    ( DownstreamStackBusLane[60][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane10_strm0_ready         ( DownstreamStackBusLane[60][10].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane10_strm0_cntl          ( DownstreamStackBusLane[60][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane10_strm0_data          ( DownstreamStackBusLane[60][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane10_strm0_data_valid    ( DownstreamStackBusLane[60][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane10_strm1_ready         ( DownstreamStackBusLane[60][10].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane10_strm1_cntl          ( DownstreamStackBusLane[60][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane10_strm1_data          ( DownstreamStackBusLane[60][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane10_strm1_data_valid    ( DownstreamStackBusLane[60][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane11_strm0_ready         ( DownstreamStackBusLane[60][11].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane11_strm0_cntl          ( DownstreamStackBusLane[60][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane11_strm0_data          ( DownstreamStackBusLane[60][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane11_strm0_data_valid    ( DownstreamStackBusLane[60][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane11_strm1_ready         ( DownstreamStackBusLane[60][11].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane11_strm1_cntl          ( DownstreamStackBusLane[60][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane11_strm1_data          ( DownstreamStackBusLane[60][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane11_strm1_data_valid    ( DownstreamStackBusLane[60][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane12_strm0_ready         ( DownstreamStackBusLane[60][12].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane12_strm0_cntl          ( DownstreamStackBusLane[60][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane12_strm0_data          ( DownstreamStackBusLane[60][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane12_strm0_data_valid    ( DownstreamStackBusLane[60][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane12_strm1_ready         ( DownstreamStackBusLane[60][12].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane12_strm1_cntl          ( DownstreamStackBusLane[60][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane12_strm1_data          ( DownstreamStackBusLane[60][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane12_strm1_data_valid    ( DownstreamStackBusLane[60][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane13_strm0_ready         ( DownstreamStackBusLane[60][13].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane13_strm0_cntl          ( DownstreamStackBusLane[60][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane13_strm0_data          ( DownstreamStackBusLane[60][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane13_strm0_data_valid    ( DownstreamStackBusLane[60][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane13_strm1_ready         ( DownstreamStackBusLane[60][13].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane13_strm1_cntl          ( DownstreamStackBusLane[60][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane13_strm1_data          ( DownstreamStackBusLane[60][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane13_strm1_data_valid    ( DownstreamStackBusLane[60][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane14_strm0_ready         ( DownstreamStackBusLane[60][14].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane14_strm0_cntl          ( DownstreamStackBusLane[60][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane14_strm0_data          ( DownstreamStackBusLane[60][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane14_strm0_data_valid    ( DownstreamStackBusLane[60][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane14_strm1_ready         ( DownstreamStackBusLane[60][14].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane14_strm1_cntl          ( DownstreamStackBusLane[60][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane14_strm1_data          ( DownstreamStackBusLane[60][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane14_strm1_data_valid    ( DownstreamStackBusLane[60][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane15_strm0_ready         ( DownstreamStackBusLane[60][15].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane15_strm0_cntl          ( DownstreamStackBusLane[60][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane15_strm0_data          ( DownstreamStackBusLane[60][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane15_strm0_data_valid    ( DownstreamStackBusLane[60][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane15_strm1_ready         ( DownstreamStackBusLane[60][15].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane15_strm1_cntl          ( DownstreamStackBusLane[60][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane15_strm1_data          ( DownstreamStackBusLane[60][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane15_strm1_data_valid    ( DownstreamStackBusLane[60][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane16_strm0_ready         ( DownstreamStackBusLane[60][16].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane16_strm0_cntl          ( DownstreamStackBusLane[60][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane16_strm0_data          ( DownstreamStackBusLane[60][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane16_strm0_data_valid    ( DownstreamStackBusLane[60][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane16_strm1_ready         ( DownstreamStackBusLane[60][16].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane16_strm1_cntl          ( DownstreamStackBusLane[60][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane16_strm1_data          ( DownstreamStackBusLane[60][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane16_strm1_data_valid    ( DownstreamStackBusLane[60][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane17_strm0_ready         ( DownstreamStackBusLane[60][17].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane17_strm0_cntl          ( DownstreamStackBusLane[60][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane17_strm0_data          ( DownstreamStackBusLane[60][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane17_strm0_data_valid    ( DownstreamStackBusLane[60][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane17_strm1_ready         ( DownstreamStackBusLane[60][17].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane17_strm1_cntl          ( DownstreamStackBusLane[60][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane17_strm1_data          ( DownstreamStackBusLane[60][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane17_strm1_data_valid    ( DownstreamStackBusLane[60][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane18_strm0_ready         ( DownstreamStackBusLane[60][18].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane18_strm0_cntl          ( DownstreamStackBusLane[60][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane18_strm0_data          ( DownstreamStackBusLane[60][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane18_strm0_data_valid    ( DownstreamStackBusLane[60][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane18_strm1_ready         ( DownstreamStackBusLane[60][18].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane18_strm1_cntl          ( DownstreamStackBusLane[60][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane18_strm1_data          ( DownstreamStackBusLane[60][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane18_strm1_data_valid    ( DownstreamStackBusLane[60][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane19_strm0_ready         ( DownstreamStackBusLane[60][19].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane19_strm0_cntl          ( DownstreamStackBusLane[60][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane19_strm0_data          ( DownstreamStackBusLane[60][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane19_strm0_data_valid    ( DownstreamStackBusLane[60][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane19_strm1_ready         ( DownstreamStackBusLane[60][19].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane19_strm1_cntl          ( DownstreamStackBusLane[60][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane19_strm1_data          ( DownstreamStackBusLane[60][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane19_strm1_data_valid    ( DownstreamStackBusLane[60][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane20_strm0_ready         ( DownstreamStackBusLane[60][20].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane20_strm0_cntl          ( DownstreamStackBusLane[60][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane20_strm0_data          ( DownstreamStackBusLane[60][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane20_strm0_data_valid    ( DownstreamStackBusLane[60][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane20_strm1_ready         ( DownstreamStackBusLane[60][20].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane20_strm1_cntl          ( DownstreamStackBusLane[60][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane20_strm1_data          ( DownstreamStackBusLane[60][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane20_strm1_data_valid    ( DownstreamStackBusLane[60][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane21_strm0_ready         ( DownstreamStackBusLane[60][21].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane21_strm0_cntl          ( DownstreamStackBusLane[60][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane21_strm0_data          ( DownstreamStackBusLane[60][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane21_strm0_data_valid    ( DownstreamStackBusLane[60][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane21_strm1_ready         ( DownstreamStackBusLane[60][21].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane21_strm1_cntl          ( DownstreamStackBusLane[60][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane21_strm1_data          ( DownstreamStackBusLane[60][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane21_strm1_data_valid    ( DownstreamStackBusLane[60][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane22_strm0_ready         ( DownstreamStackBusLane[60][22].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane22_strm0_cntl          ( DownstreamStackBusLane[60][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane22_strm0_data          ( DownstreamStackBusLane[60][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane22_strm0_data_valid    ( DownstreamStackBusLane[60][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane22_strm1_ready         ( DownstreamStackBusLane[60][22].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane22_strm1_cntl          ( DownstreamStackBusLane[60][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane22_strm1_data          ( DownstreamStackBusLane[60][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane22_strm1_data_valid    ( DownstreamStackBusLane[60][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane23_strm0_ready         ( DownstreamStackBusLane[60][23].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane23_strm0_cntl          ( DownstreamStackBusLane[60][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane23_strm0_data          ( DownstreamStackBusLane[60][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane23_strm0_data_valid    ( DownstreamStackBusLane[60][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane23_strm1_ready         ( DownstreamStackBusLane[60][23].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane23_strm1_cntl          ( DownstreamStackBusLane[60][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane23_strm1_data          ( DownstreamStackBusLane[60][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane23_strm1_data_valid    ( DownstreamStackBusLane[60][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane24_strm0_ready         ( DownstreamStackBusLane[60][24].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane24_strm0_cntl          ( DownstreamStackBusLane[60][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane24_strm0_data          ( DownstreamStackBusLane[60][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane24_strm0_data_valid    ( DownstreamStackBusLane[60][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane24_strm1_ready         ( DownstreamStackBusLane[60][24].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane24_strm1_cntl          ( DownstreamStackBusLane[60][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane24_strm1_data          ( DownstreamStackBusLane[60][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane24_strm1_data_valid    ( DownstreamStackBusLane[60][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane25_strm0_ready         ( DownstreamStackBusLane[60][25].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane25_strm0_cntl          ( DownstreamStackBusLane[60][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane25_strm0_data          ( DownstreamStackBusLane[60][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane25_strm0_data_valid    ( DownstreamStackBusLane[60][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane25_strm1_ready         ( DownstreamStackBusLane[60][25].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane25_strm1_cntl          ( DownstreamStackBusLane[60][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane25_strm1_data          ( DownstreamStackBusLane[60][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane25_strm1_data_valid    ( DownstreamStackBusLane[60][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane26_strm0_ready         ( DownstreamStackBusLane[60][26].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane26_strm0_cntl          ( DownstreamStackBusLane[60][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane26_strm0_data          ( DownstreamStackBusLane[60][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane26_strm0_data_valid    ( DownstreamStackBusLane[60][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane26_strm1_ready         ( DownstreamStackBusLane[60][26].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane26_strm1_cntl          ( DownstreamStackBusLane[60][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane26_strm1_data          ( DownstreamStackBusLane[60][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane26_strm1_data_valid    ( DownstreamStackBusLane[60][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane27_strm0_ready         ( DownstreamStackBusLane[60][27].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane27_strm0_cntl          ( DownstreamStackBusLane[60][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane27_strm0_data          ( DownstreamStackBusLane[60][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane27_strm0_data_valid    ( DownstreamStackBusLane[60][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane27_strm1_ready         ( DownstreamStackBusLane[60][27].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane27_strm1_cntl          ( DownstreamStackBusLane[60][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane27_strm1_data          ( DownstreamStackBusLane[60][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane27_strm1_data_valid    ( DownstreamStackBusLane[60][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane28_strm0_ready         ( DownstreamStackBusLane[60][28].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane28_strm0_cntl          ( DownstreamStackBusLane[60][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane28_strm0_data          ( DownstreamStackBusLane[60][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane28_strm0_data_valid    ( DownstreamStackBusLane[60][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane28_strm1_ready         ( DownstreamStackBusLane[60][28].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane28_strm1_cntl          ( DownstreamStackBusLane[60][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane28_strm1_data          ( DownstreamStackBusLane[60][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane28_strm1_data_valid    ( DownstreamStackBusLane[60][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane29_strm0_ready         ( DownstreamStackBusLane[60][29].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane29_strm0_cntl          ( DownstreamStackBusLane[60][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane29_strm0_data          ( DownstreamStackBusLane[60][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane29_strm0_data_valid    ( DownstreamStackBusLane[60][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane29_strm1_ready         ( DownstreamStackBusLane[60][29].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane29_strm1_cntl          ( DownstreamStackBusLane[60][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane29_strm1_data          ( DownstreamStackBusLane[60][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane29_strm1_data_valid    ( DownstreamStackBusLane[60][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane30_strm0_ready         ( DownstreamStackBusLane[60][30].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane30_strm0_cntl          ( DownstreamStackBusLane[60][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane30_strm0_data          ( DownstreamStackBusLane[60][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane30_strm0_data_valid    ( DownstreamStackBusLane[60][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane30_strm1_ready         ( DownstreamStackBusLane[60][30].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane30_strm1_cntl          ( DownstreamStackBusLane[60][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane30_strm1_data          ( DownstreamStackBusLane[60][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane30_strm1_data_valid    ( DownstreamStackBusLane[60][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 60, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane31_strm0_ready         ( DownstreamStackBusLane[60][31].pe__std__lane_strm0_ready              ),      
        .std__pe60__lane31_strm0_cntl          ( DownstreamStackBusLane[60][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe60__lane31_strm0_data          ( DownstreamStackBusLane[60][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe60__lane31_strm0_data_valid    ( DownstreamStackBusLane[60][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__std__lane31_strm1_ready         ( DownstreamStackBusLane[60][31].pe__std__lane_strm1_ready              ),      
        .std__pe60__lane31_strm1_cntl          ( DownstreamStackBusLane[60][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe60__lane31_strm1_data          ( DownstreamStackBusLane[60][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe60__lane31_strm1_data_valid    ( DownstreamStackBusLane[60][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane0_strm0_ready         ( DownstreamStackBusLane[61][0].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane0_strm0_cntl          ( DownstreamStackBusLane[61][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane0_strm0_data          ( DownstreamStackBusLane[61][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane0_strm0_data_valid    ( DownstreamStackBusLane[61][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane0_strm1_ready         ( DownstreamStackBusLane[61][0].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane0_strm1_cntl          ( DownstreamStackBusLane[61][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane0_strm1_data          ( DownstreamStackBusLane[61][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane0_strm1_data_valid    ( DownstreamStackBusLane[61][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane1_strm0_ready         ( DownstreamStackBusLane[61][1].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane1_strm0_cntl          ( DownstreamStackBusLane[61][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane1_strm0_data          ( DownstreamStackBusLane[61][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane1_strm0_data_valid    ( DownstreamStackBusLane[61][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane1_strm1_ready         ( DownstreamStackBusLane[61][1].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane1_strm1_cntl          ( DownstreamStackBusLane[61][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane1_strm1_data          ( DownstreamStackBusLane[61][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane1_strm1_data_valid    ( DownstreamStackBusLane[61][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane2_strm0_ready         ( DownstreamStackBusLane[61][2].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane2_strm0_cntl          ( DownstreamStackBusLane[61][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane2_strm0_data          ( DownstreamStackBusLane[61][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane2_strm0_data_valid    ( DownstreamStackBusLane[61][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane2_strm1_ready         ( DownstreamStackBusLane[61][2].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane2_strm1_cntl          ( DownstreamStackBusLane[61][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane2_strm1_data          ( DownstreamStackBusLane[61][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane2_strm1_data_valid    ( DownstreamStackBusLane[61][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane3_strm0_ready         ( DownstreamStackBusLane[61][3].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane3_strm0_cntl          ( DownstreamStackBusLane[61][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane3_strm0_data          ( DownstreamStackBusLane[61][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane3_strm0_data_valid    ( DownstreamStackBusLane[61][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane3_strm1_ready         ( DownstreamStackBusLane[61][3].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane3_strm1_cntl          ( DownstreamStackBusLane[61][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane3_strm1_data          ( DownstreamStackBusLane[61][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane3_strm1_data_valid    ( DownstreamStackBusLane[61][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane4_strm0_ready         ( DownstreamStackBusLane[61][4].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane4_strm0_cntl          ( DownstreamStackBusLane[61][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane4_strm0_data          ( DownstreamStackBusLane[61][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane4_strm0_data_valid    ( DownstreamStackBusLane[61][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane4_strm1_ready         ( DownstreamStackBusLane[61][4].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane4_strm1_cntl          ( DownstreamStackBusLane[61][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane4_strm1_data          ( DownstreamStackBusLane[61][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane4_strm1_data_valid    ( DownstreamStackBusLane[61][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane5_strm0_ready         ( DownstreamStackBusLane[61][5].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane5_strm0_cntl          ( DownstreamStackBusLane[61][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane5_strm0_data          ( DownstreamStackBusLane[61][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane5_strm0_data_valid    ( DownstreamStackBusLane[61][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane5_strm1_ready         ( DownstreamStackBusLane[61][5].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane5_strm1_cntl          ( DownstreamStackBusLane[61][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane5_strm1_data          ( DownstreamStackBusLane[61][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane5_strm1_data_valid    ( DownstreamStackBusLane[61][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane6_strm0_ready         ( DownstreamStackBusLane[61][6].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane6_strm0_cntl          ( DownstreamStackBusLane[61][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane6_strm0_data          ( DownstreamStackBusLane[61][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane6_strm0_data_valid    ( DownstreamStackBusLane[61][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane6_strm1_ready         ( DownstreamStackBusLane[61][6].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane6_strm1_cntl          ( DownstreamStackBusLane[61][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane6_strm1_data          ( DownstreamStackBusLane[61][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane6_strm1_data_valid    ( DownstreamStackBusLane[61][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane7_strm0_ready         ( DownstreamStackBusLane[61][7].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane7_strm0_cntl          ( DownstreamStackBusLane[61][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane7_strm0_data          ( DownstreamStackBusLane[61][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane7_strm0_data_valid    ( DownstreamStackBusLane[61][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane7_strm1_ready         ( DownstreamStackBusLane[61][7].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane7_strm1_cntl          ( DownstreamStackBusLane[61][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane7_strm1_data          ( DownstreamStackBusLane[61][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane7_strm1_data_valid    ( DownstreamStackBusLane[61][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane8_strm0_ready         ( DownstreamStackBusLane[61][8].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane8_strm0_cntl          ( DownstreamStackBusLane[61][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane8_strm0_data          ( DownstreamStackBusLane[61][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane8_strm0_data_valid    ( DownstreamStackBusLane[61][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane8_strm1_ready         ( DownstreamStackBusLane[61][8].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane8_strm1_cntl          ( DownstreamStackBusLane[61][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane8_strm1_data          ( DownstreamStackBusLane[61][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane8_strm1_data_valid    ( DownstreamStackBusLane[61][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane9_strm0_ready         ( DownstreamStackBusLane[61][9].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane9_strm0_cntl          ( DownstreamStackBusLane[61][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane9_strm0_data          ( DownstreamStackBusLane[61][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane9_strm0_data_valid    ( DownstreamStackBusLane[61][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane9_strm1_ready         ( DownstreamStackBusLane[61][9].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane9_strm1_cntl          ( DownstreamStackBusLane[61][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane9_strm1_data          ( DownstreamStackBusLane[61][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane9_strm1_data_valid    ( DownstreamStackBusLane[61][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane10_strm0_ready         ( DownstreamStackBusLane[61][10].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane10_strm0_cntl          ( DownstreamStackBusLane[61][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane10_strm0_data          ( DownstreamStackBusLane[61][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane10_strm0_data_valid    ( DownstreamStackBusLane[61][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane10_strm1_ready         ( DownstreamStackBusLane[61][10].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane10_strm1_cntl          ( DownstreamStackBusLane[61][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane10_strm1_data          ( DownstreamStackBusLane[61][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane10_strm1_data_valid    ( DownstreamStackBusLane[61][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane11_strm0_ready         ( DownstreamStackBusLane[61][11].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane11_strm0_cntl          ( DownstreamStackBusLane[61][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane11_strm0_data          ( DownstreamStackBusLane[61][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane11_strm0_data_valid    ( DownstreamStackBusLane[61][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane11_strm1_ready         ( DownstreamStackBusLane[61][11].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane11_strm1_cntl          ( DownstreamStackBusLane[61][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane11_strm1_data          ( DownstreamStackBusLane[61][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane11_strm1_data_valid    ( DownstreamStackBusLane[61][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane12_strm0_ready         ( DownstreamStackBusLane[61][12].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane12_strm0_cntl          ( DownstreamStackBusLane[61][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane12_strm0_data          ( DownstreamStackBusLane[61][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane12_strm0_data_valid    ( DownstreamStackBusLane[61][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane12_strm1_ready         ( DownstreamStackBusLane[61][12].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane12_strm1_cntl          ( DownstreamStackBusLane[61][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane12_strm1_data          ( DownstreamStackBusLane[61][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane12_strm1_data_valid    ( DownstreamStackBusLane[61][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane13_strm0_ready         ( DownstreamStackBusLane[61][13].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane13_strm0_cntl          ( DownstreamStackBusLane[61][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane13_strm0_data          ( DownstreamStackBusLane[61][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane13_strm0_data_valid    ( DownstreamStackBusLane[61][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane13_strm1_ready         ( DownstreamStackBusLane[61][13].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane13_strm1_cntl          ( DownstreamStackBusLane[61][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane13_strm1_data          ( DownstreamStackBusLane[61][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane13_strm1_data_valid    ( DownstreamStackBusLane[61][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane14_strm0_ready         ( DownstreamStackBusLane[61][14].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane14_strm0_cntl          ( DownstreamStackBusLane[61][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane14_strm0_data          ( DownstreamStackBusLane[61][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane14_strm0_data_valid    ( DownstreamStackBusLane[61][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane14_strm1_ready         ( DownstreamStackBusLane[61][14].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane14_strm1_cntl          ( DownstreamStackBusLane[61][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane14_strm1_data          ( DownstreamStackBusLane[61][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane14_strm1_data_valid    ( DownstreamStackBusLane[61][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane15_strm0_ready         ( DownstreamStackBusLane[61][15].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane15_strm0_cntl          ( DownstreamStackBusLane[61][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane15_strm0_data          ( DownstreamStackBusLane[61][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane15_strm0_data_valid    ( DownstreamStackBusLane[61][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane15_strm1_ready         ( DownstreamStackBusLane[61][15].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane15_strm1_cntl          ( DownstreamStackBusLane[61][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane15_strm1_data          ( DownstreamStackBusLane[61][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane15_strm1_data_valid    ( DownstreamStackBusLane[61][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane16_strm0_ready         ( DownstreamStackBusLane[61][16].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane16_strm0_cntl          ( DownstreamStackBusLane[61][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane16_strm0_data          ( DownstreamStackBusLane[61][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane16_strm0_data_valid    ( DownstreamStackBusLane[61][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane16_strm1_ready         ( DownstreamStackBusLane[61][16].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane16_strm1_cntl          ( DownstreamStackBusLane[61][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane16_strm1_data          ( DownstreamStackBusLane[61][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane16_strm1_data_valid    ( DownstreamStackBusLane[61][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane17_strm0_ready         ( DownstreamStackBusLane[61][17].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane17_strm0_cntl          ( DownstreamStackBusLane[61][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane17_strm0_data          ( DownstreamStackBusLane[61][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane17_strm0_data_valid    ( DownstreamStackBusLane[61][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane17_strm1_ready         ( DownstreamStackBusLane[61][17].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane17_strm1_cntl          ( DownstreamStackBusLane[61][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane17_strm1_data          ( DownstreamStackBusLane[61][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane17_strm1_data_valid    ( DownstreamStackBusLane[61][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane18_strm0_ready         ( DownstreamStackBusLane[61][18].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane18_strm0_cntl          ( DownstreamStackBusLane[61][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane18_strm0_data          ( DownstreamStackBusLane[61][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane18_strm0_data_valid    ( DownstreamStackBusLane[61][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane18_strm1_ready         ( DownstreamStackBusLane[61][18].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane18_strm1_cntl          ( DownstreamStackBusLane[61][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane18_strm1_data          ( DownstreamStackBusLane[61][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane18_strm1_data_valid    ( DownstreamStackBusLane[61][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane19_strm0_ready         ( DownstreamStackBusLane[61][19].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane19_strm0_cntl          ( DownstreamStackBusLane[61][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane19_strm0_data          ( DownstreamStackBusLane[61][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane19_strm0_data_valid    ( DownstreamStackBusLane[61][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane19_strm1_ready         ( DownstreamStackBusLane[61][19].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane19_strm1_cntl          ( DownstreamStackBusLane[61][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane19_strm1_data          ( DownstreamStackBusLane[61][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane19_strm1_data_valid    ( DownstreamStackBusLane[61][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane20_strm0_ready         ( DownstreamStackBusLane[61][20].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane20_strm0_cntl          ( DownstreamStackBusLane[61][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane20_strm0_data          ( DownstreamStackBusLane[61][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane20_strm0_data_valid    ( DownstreamStackBusLane[61][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane20_strm1_ready         ( DownstreamStackBusLane[61][20].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane20_strm1_cntl          ( DownstreamStackBusLane[61][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane20_strm1_data          ( DownstreamStackBusLane[61][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane20_strm1_data_valid    ( DownstreamStackBusLane[61][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane21_strm0_ready         ( DownstreamStackBusLane[61][21].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane21_strm0_cntl          ( DownstreamStackBusLane[61][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane21_strm0_data          ( DownstreamStackBusLane[61][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane21_strm0_data_valid    ( DownstreamStackBusLane[61][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane21_strm1_ready         ( DownstreamStackBusLane[61][21].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane21_strm1_cntl          ( DownstreamStackBusLane[61][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane21_strm1_data          ( DownstreamStackBusLane[61][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane21_strm1_data_valid    ( DownstreamStackBusLane[61][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane22_strm0_ready         ( DownstreamStackBusLane[61][22].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane22_strm0_cntl          ( DownstreamStackBusLane[61][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane22_strm0_data          ( DownstreamStackBusLane[61][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane22_strm0_data_valid    ( DownstreamStackBusLane[61][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane22_strm1_ready         ( DownstreamStackBusLane[61][22].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane22_strm1_cntl          ( DownstreamStackBusLane[61][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane22_strm1_data          ( DownstreamStackBusLane[61][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane22_strm1_data_valid    ( DownstreamStackBusLane[61][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane23_strm0_ready         ( DownstreamStackBusLane[61][23].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane23_strm0_cntl          ( DownstreamStackBusLane[61][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane23_strm0_data          ( DownstreamStackBusLane[61][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane23_strm0_data_valid    ( DownstreamStackBusLane[61][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane23_strm1_ready         ( DownstreamStackBusLane[61][23].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane23_strm1_cntl          ( DownstreamStackBusLane[61][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane23_strm1_data          ( DownstreamStackBusLane[61][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane23_strm1_data_valid    ( DownstreamStackBusLane[61][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane24_strm0_ready         ( DownstreamStackBusLane[61][24].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane24_strm0_cntl          ( DownstreamStackBusLane[61][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane24_strm0_data          ( DownstreamStackBusLane[61][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane24_strm0_data_valid    ( DownstreamStackBusLane[61][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane24_strm1_ready         ( DownstreamStackBusLane[61][24].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane24_strm1_cntl          ( DownstreamStackBusLane[61][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane24_strm1_data          ( DownstreamStackBusLane[61][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane24_strm1_data_valid    ( DownstreamStackBusLane[61][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane25_strm0_ready         ( DownstreamStackBusLane[61][25].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane25_strm0_cntl          ( DownstreamStackBusLane[61][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane25_strm0_data          ( DownstreamStackBusLane[61][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane25_strm0_data_valid    ( DownstreamStackBusLane[61][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane25_strm1_ready         ( DownstreamStackBusLane[61][25].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane25_strm1_cntl          ( DownstreamStackBusLane[61][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane25_strm1_data          ( DownstreamStackBusLane[61][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane25_strm1_data_valid    ( DownstreamStackBusLane[61][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane26_strm0_ready         ( DownstreamStackBusLane[61][26].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane26_strm0_cntl          ( DownstreamStackBusLane[61][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane26_strm0_data          ( DownstreamStackBusLane[61][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane26_strm0_data_valid    ( DownstreamStackBusLane[61][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane26_strm1_ready         ( DownstreamStackBusLane[61][26].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane26_strm1_cntl          ( DownstreamStackBusLane[61][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane26_strm1_data          ( DownstreamStackBusLane[61][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane26_strm1_data_valid    ( DownstreamStackBusLane[61][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane27_strm0_ready         ( DownstreamStackBusLane[61][27].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane27_strm0_cntl          ( DownstreamStackBusLane[61][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane27_strm0_data          ( DownstreamStackBusLane[61][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane27_strm0_data_valid    ( DownstreamStackBusLane[61][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane27_strm1_ready         ( DownstreamStackBusLane[61][27].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane27_strm1_cntl          ( DownstreamStackBusLane[61][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane27_strm1_data          ( DownstreamStackBusLane[61][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane27_strm1_data_valid    ( DownstreamStackBusLane[61][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane28_strm0_ready         ( DownstreamStackBusLane[61][28].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane28_strm0_cntl          ( DownstreamStackBusLane[61][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane28_strm0_data          ( DownstreamStackBusLane[61][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane28_strm0_data_valid    ( DownstreamStackBusLane[61][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane28_strm1_ready         ( DownstreamStackBusLane[61][28].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane28_strm1_cntl          ( DownstreamStackBusLane[61][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane28_strm1_data          ( DownstreamStackBusLane[61][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane28_strm1_data_valid    ( DownstreamStackBusLane[61][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane29_strm0_ready         ( DownstreamStackBusLane[61][29].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane29_strm0_cntl          ( DownstreamStackBusLane[61][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane29_strm0_data          ( DownstreamStackBusLane[61][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane29_strm0_data_valid    ( DownstreamStackBusLane[61][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane29_strm1_ready         ( DownstreamStackBusLane[61][29].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane29_strm1_cntl          ( DownstreamStackBusLane[61][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane29_strm1_data          ( DownstreamStackBusLane[61][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane29_strm1_data_valid    ( DownstreamStackBusLane[61][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane30_strm0_ready         ( DownstreamStackBusLane[61][30].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane30_strm0_cntl          ( DownstreamStackBusLane[61][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane30_strm0_data          ( DownstreamStackBusLane[61][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane30_strm0_data_valid    ( DownstreamStackBusLane[61][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane30_strm1_ready         ( DownstreamStackBusLane[61][30].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane30_strm1_cntl          ( DownstreamStackBusLane[61][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane30_strm1_data          ( DownstreamStackBusLane[61][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane30_strm1_data_valid    ( DownstreamStackBusLane[61][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 61, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane31_strm0_ready         ( DownstreamStackBusLane[61][31].pe__std__lane_strm0_ready              ),      
        .std__pe61__lane31_strm0_cntl          ( DownstreamStackBusLane[61][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe61__lane31_strm0_data          ( DownstreamStackBusLane[61][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe61__lane31_strm0_data_valid    ( DownstreamStackBusLane[61][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__std__lane31_strm1_ready         ( DownstreamStackBusLane[61][31].pe__std__lane_strm1_ready              ),      
        .std__pe61__lane31_strm1_cntl          ( DownstreamStackBusLane[61][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe61__lane31_strm1_data          ( DownstreamStackBusLane[61][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe61__lane31_strm1_data_valid    ( DownstreamStackBusLane[61][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane0_strm0_ready         ( DownstreamStackBusLane[62][0].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane0_strm0_cntl          ( DownstreamStackBusLane[62][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane0_strm0_data          ( DownstreamStackBusLane[62][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane0_strm0_data_valid    ( DownstreamStackBusLane[62][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane0_strm1_ready         ( DownstreamStackBusLane[62][0].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane0_strm1_cntl          ( DownstreamStackBusLane[62][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane0_strm1_data          ( DownstreamStackBusLane[62][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane0_strm1_data_valid    ( DownstreamStackBusLane[62][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane1_strm0_ready         ( DownstreamStackBusLane[62][1].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane1_strm0_cntl          ( DownstreamStackBusLane[62][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane1_strm0_data          ( DownstreamStackBusLane[62][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane1_strm0_data_valid    ( DownstreamStackBusLane[62][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane1_strm1_ready         ( DownstreamStackBusLane[62][1].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane1_strm1_cntl          ( DownstreamStackBusLane[62][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane1_strm1_data          ( DownstreamStackBusLane[62][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane1_strm1_data_valid    ( DownstreamStackBusLane[62][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane2_strm0_ready         ( DownstreamStackBusLane[62][2].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane2_strm0_cntl          ( DownstreamStackBusLane[62][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane2_strm0_data          ( DownstreamStackBusLane[62][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane2_strm0_data_valid    ( DownstreamStackBusLane[62][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane2_strm1_ready         ( DownstreamStackBusLane[62][2].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane2_strm1_cntl          ( DownstreamStackBusLane[62][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane2_strm1_data          ( DownstreamStackBusLane[62][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane2_strm1_data_valid    ( DownstreamStackBusLane[62][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane3_strm0_ready         ( DownstreamStackBusLane[62][3].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane3_strm0_cntl          ( DownstreamStackBusLane[62][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane3_strm0_data          ( DownstreamStackBusLane[62][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane3_strm0_data_valid    ( DownstreamStackBusLane[62][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane3_strm1_ready         ( DownstreamStackBusLane[62][3].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane3_strm1_cntl          ( DownstreamStackBusLane[62][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane3_strm1_data          ( DownstreamStackBusLane[62][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane3_strm1_data_valid    ( DownstreamStackBusLane[62][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane4_strm0_ready         ( DownstreamStackBusLane[62][4].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane4_strm0_cntl          ( DownstreamStackBusLane[62][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane4_strm0_data          ( DownstreamStackBusLane[62][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane4_strm0_data_valid    ( DownstreamStackBusLane[62][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane4_strm1_ready         ( DownstreamStackBusLane[62][4].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane4_strm1_cntl          ( DownstreamStackBusLane[62][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane4_strm1_data          ( DownstreamStackBusLane[62][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane4_strm1_data_valid    ( DownstreamStackBusLane[62][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane5_strm0_ready         ( DownstreamStackBusLane[62][5].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane5_strm0_cntl          ( DownstreamStackBusLane[62][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane5_strm0_data          ( DownstreamStackBusLane[62][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane5_strm0_data_valid    ( DownstreamStackBusLane[62][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane5_strm1_ready         ( DownstreamStackBusLane[62][5].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane5_strm1_cntl          ( DownstreamStackBusLane[62][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane5_strm1_data          ( DownstreamStackBusLane[62][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane5_strm1_data_valid    ( DownstreamStackBusLane[62][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane6_strm0_ready         ( DownstreamStackBusLane[62][6].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane6_strm0_cntl          ( DownstreamStackBusLane[62][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane6_strm0_data          ( DownstreamStackBusLane[62][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane6_strm0_data_valid    ( DownstreamStackBusLane[62][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane6_strm1_ready         ( DownstreamStackBusLane[62][6].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane6_strm1_cntl          ( DownstreamStackBusLane[62][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane6_strm1_data          ( DownstreamStackBusLane[62][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane6_strm1_data_valid    ( DownstreamStackBusLane[62][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane7_strm0_ready         ( DownstreamStackBusLane[62][7].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane7_strm0_cntl          ( DownstreamStackBusLane[62][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane7_strm0_data          ( DownstreamStackBusLane[62][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane7_strm0_data_valid    ( DownstreamStackBusLane[62][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane7_strm1_ready         ( DownstreamStackBusLane[62][7].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane7_strm1_cntl          ( DownstreamStackBusLane[62][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane7_strm1_data          ( DownstreamStackBusLane[62][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane7_strm1_data_valid    ( DownstreamStackBusLane[62][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane8_strm0_ready         ( DownstreamStackBusLane[62][8].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane8_strm0_cntl          ( DownstreamStackBusLane[62][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane8_strm0_data          ( DownstreamStackBusLane[62][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane8_strm0_data_valid    ( DownstreamStackBusLane[62][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane8_strm1_ready         ( DownstreamStackBusLane[62][8].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane8_strm1_cntl          ( DownstreamStackBusLane[62][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane8_strm1_data          ( DownstreamStackBusLane[62][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane8_strm1_data_valid    ( DownstreamStackBusLane[62][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane9_strm0_ready         ( DownstreamStackBusLane[62][9].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane9_strm0_cntl          ( DownstreamStackBusLane[62][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane9_strm0_data          ( DownstreamStackBusLane[62][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane9_strm0_data_valid    ( DownstreamStackBusLane[62][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane9_strm1_ready         ( DownstreamStackBusLane[62][9].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane9_strm1_cntl          ( DownstreamStackBusLane[62][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane9_strm1_data          ( DownstreamStackBusLane[62][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane9_strm1_data_valid    ( DownstreamStackBusLane[62][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane10_strm0_ready         ( DownstreamStackBusLane[62][10].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane10_strm0_cntl          ( DownstreamStackBusLane[62][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane10_strm0_data          ( DownstreamStackBusLane[62][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane10_strm0_data_valid    ( DownstreamStackBusLane[62][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane10_strm1_ready         ( DownstreamStackBusLane[62][10].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane10_strm1_cntl          ( DownstreamStackBusLane[62][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane10_strm1_data          ( DownstreamStackBusLane[62][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane10_strm1_data_valid    ( DownstreamStackBusLane[62][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane11_strm0_ready         ( DownstreamStackBusLane[62][11].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane11_strm0_cntl          ( DownstreamStackBusLane[62][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane11_strm0_data          ( DownstreamStackBusLane[62][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane11_strm0_data_valid    ( DownstreamStackBusLane[62][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane11_strm1_ready         ( DownstreamStackBusLane[62][11].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane11_strm1_cntl          ( DownstreamStackBusLane[62][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane11_strm1_data          ( DownstreamStackBusLane[62][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane11_strm1_data_valid    ( DownstreamStackBusLane[62][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane12_strm0_ready         ( DownstreamStackBusLane[62][12].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane12_strm0_cntl          ( DownstreamStackBusLane[62][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane12_strm0_data          ( DownstreamStackBusLane[62][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane12_strm0_data_valid    ( DownstreamStackBusLane[62][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane12_strm1_ready         ( DownstreamStackBusLane[62][12].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane12_strm1_cntl          ( DownstreamStackBusLane[62][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane12_strm1_data          ( DownstreamStackBusLane[62][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane12_strm1_data_valid    ( DownstreamStackBusLane[62][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane13_strm0_ready         ( DownstreamStackBusLane[62][13].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane13_strm0_cntl          ( DownstreamStackBusLane[62][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane13_strm0_data          ( DownstreamStackBusLane[62][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane13_strm0_data_valid    ( DownstreamStackBusLane[62][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane13_strm1_ready         ( DownstreamStackBusLane[62][13].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane13_strm1_cntl          ( DownstreamStackBusLane[62][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane13_strm1_data          ( DownstreamStackBusLane[62][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane13_strm1_data_valid    ( DownstreamStackBusLane[62][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane14_strm0_ready         ( DownstreamStackBusLane[62][14].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane14_strm0_cntl          ( DownstreamStackBusLane[62][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane14_strm0_data          ( DownstreamStackBusLane[62][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane14_strm0_data_valid    ( DownstreamStackBusLane[62][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane14_strm1_ready         ( DownstreamStackBusLane[62][14].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane14_strm1_cntl          ( DownstreamStackBusLane[62][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane14_strm1_data          ( DownstreamStackBusLane[62][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane14_strm1_data_valid    ( DownstreamStackBusLane[62][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane15_strm0_ready         ( DownstreamStackBusLane[62][15].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane15_strm0_cntl          ( DownstreamStackBusLane[62][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane15_strm0_data          ( DownstreamStackBusLane[62][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane15_strm0_data_valid    ( DownstreamStackBusLane[62][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane15_strm1_ready         ( DownstreamStackBusLane[62][15].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane15_strm1_cntl          ( DownstreamStackBusLane[62][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane15_strm1_data          ( DownstreamStackBusLane[62][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane15_strm1_data_valid    ( DownstreamStackBusLane[62][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane16_strm0_ready         ( DownstreamStackBusLane[62][16].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane16_strm0_cntl          ( DownstreamStackBusLane[62][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane16_strm0_data          ( DownstreamStackBusLane[62][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane16_strm0_data_valid    ( DownstreamStackBusLane[62][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane16_strm1_ready         ( DownstreamStackBusLane[62][16].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane16_strm1_cntl          ( DownstreamStackBusLane[62][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane16_strm1_data          ( DownstreamStackBusLane[62][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane16_strm1_data_valid    ( DownstreamStackBusLane[62][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane17_strm0_ready         ( DownstreamStackBusLane[62][17].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane17_strm0_cntl          ( DownstreamStackBusLane[62][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane17_strm0_data          ( DownstreamStackBusLane[62][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane17_strm0_data_valid    ( DownstreamStackBusLane[62][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane17_strm1_ready         ( DownstreamStackBusLane[62][17].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane17_strm1_cntl          ( DownstreamStackBusLane[62][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane17_strm1_data          ( DownstreamStackBusLane[62][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane17_strm1_data_valid    ( DownstreamStackBusLane[62][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane18_strm0_ready         ( DownstreamStackBusLane[62][18].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane18_strm0_cntl          ( DownstreamStackBusLane[62][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane18_strm0_data          ( DownstreamStackBusLane[62][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane18_strm0_data_valid    ( DownstreamStackBusLane[62][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane18_strm1_ready         ( DownstreamStackBusLane[62][18].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane18_strm1_cntl          ( DownstreamStackBusLane[62][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane18_strm1_data          ( DownstreamStackBusLane[62][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane18_strm1_data_valid    ( DownstreamStackBusLane[62][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane19_strm0_ready         ( DownstreamStackBusLane[62][19].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane19_strm0_cntl          ( DownstreamStackBusLane[62][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane19_strm0_data          ( DownstreamStackBusLane[62][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane19_strm0_data_valid    ( DownstreamStackBusLane[62][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane19_strm1_ready         ( DownstreamStackBusLane[62][19].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane19_strm1_cntl          ( DownstreamStackBusLane[62][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane19_strm1_data          ( DownstreamStackBusLane[62][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane19_strm1_data_valid    ( DownstreamStackBusLane[62][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane20_strm0_ready         ( DownstreamStackBusLane[62][20].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane20_strm0_cntl          ( DownstreamStackBusLane[62][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane20_strm0_data          ( DownstreamStackBusLane[62][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane20_strm0_data_valid    ( DownstreamStackBusLane[62][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane20_strm1_ready         ( DownstreamStackBusLane[62][20].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane20_strm1_cntl          ( DownstreamStackBusLane[62][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane20_strm1_data          ( DownstreamStackBusLane[62][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane20_strm1_data_valid    ( DownstreamStackBusLane[62][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane21_strm0_ready         ( DownstreamStackBusLane[62][21].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane21_strm0_cntl          ( DownstreamStackBusLane[62][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane21_strm0_data          ( DownstreamStackBusLane[62][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane21_strm0_data_valid    ( DownstreamStackBusLane[62][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane21_strm1_ready         ( DownstreamStackBusLane[62][21].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane21_strm1_cntl          ( DownstreamStackBusLane[62][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane21_strm1_data          ( DownstreamStackBusLane[62][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane21_strm1_data_valid    ( DownstreamStackBusLane[62][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane22_strm0_ready         ( DownstreamStackBusLane[62][22].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane22_strm0_cntl          ( DownstreamStackBusLane[62][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane22_strm0_data          ( DownstreamStackBusLane[62][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane22_strm0_data_valid    ( DownstreamStackBusLane[62][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane22_strm1_ready         ( DownstreamStackBusLane[62][22].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane22_strm1_cntl          ( DownstreamStackBusLane[62][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane22_strm1_data          ( DownstreamStackBusLane[62][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane22_strm1_data_valid    ( DownstreamStackBusLane[62][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane23_strm0_ready         ( DownstreamStackBusLane[62][23].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane23_strm0_cntl          ( DownstreamStackBusLane[62][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane23_strm0_data          ( DownstreamStackBusLane[62][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane23_strm0_data_valid    ( DownstreamStackBusLane[62][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane23_strm1_ready         ( DownstreamStackBusLane[62][23].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane23_strm1_cntl          ( DownstreamStackBusLane[62][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane23_strm1_data          ( DownstreamStackBusLane[62][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane23_strm1_data_valid    ( DownstreamStackBusLane[62][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane24_strm0_ready         ( DownstreamStackBusLane[62][24].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane24_strm0_cntl          ( DownstreamStackBusLane[62][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane24_strm0_data          ( DownstreamStackBusLane[62][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane24_strm0_data_valid    ( DownstreamStackBusLane[62][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane24_strm1_ready         ( DownstreamStackBusLane[62][24].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane24_strm1_cntl          ( DownstreamStackBusLane[62][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane24_strm1_data          ( DownstreamStackBusLane[62][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane24_strm1_data_valid    ( DownstreamStackBusLane[62][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane25_strm0_ready         ( DownstreamStackBusLane[62][25].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane25_strm0_cntl          ( DownstreamStackBusLane[62][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane25_strm0_data          ( DownstreamStackBusLane[62][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane25_strm0_data_valid    ( DownstreamStackBusLane[62][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane25_strm1_ready         ( DownstreamStackBusLane[62][25].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane25_strm1_cntl          ( DownstreamStackBusLane[62][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane25_strm1_data          ( DownstreamStackBusLane[62][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane25_strm1_data_valid    ( DownstreamStackBusLane[62][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane26_strm0_ready         ( DownstreamStackBusLane[62][26].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane26_strm0_cntl          ( DownstreamStackBusLane[62][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane26_strm0_data          ( DownstreamStackBusLane[62][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane26_strm0_data_valid    ( DownstreamStackBusLane[62][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane26_strm1_ready         ( DownstreamStackBusLane[62][26].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane26_strm1_cntl          ( DownstreamStackBusLane[62][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane26_strm1_data          ( DownstreamStackBusLane[62][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane26_strm1_data_valid    ( DownstreamStackBusLane[62][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane27_strm0_ready         ( DownstreamStackBusLane[62][27].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane27_strm0_cntl          ( DownstreamStackBusLane[62][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane27_strm0_data          ( DownstreamStackBusLane[62][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane27_strm0_data_valid    ( DownstreamStackBusLane[62][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane27_strm1_ready         ( DownstreamStackBusLane[62][27].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane27_strm1_cntl          ( DownstreamStackBusLane[62][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane27_strm1_data          ( DownstreamStackBusLane[62][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane27_strm1_data_valid    ( DownstreamStackBusLane[62][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane28_strm0_ready         ( DownstreamStackBusLane[62][28].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane28_strm0_cntl          ( DownstreamStackBusLane[62][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane28_strm0_data          ( DownstreamStackBusLane[62][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane28_strm0_data_valid    ( DownstreamStackBusLane[62][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane28_strm1_ready         ( DownstreamStackBusLane[62][28].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane28_strm1_cntl          ( DownstreamStackBusLane[62][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane28_strm1_data          ( DownstreamStackBusLane[62][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane28_strm1_data_valid    ( DownstreamStackBusLane[62][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane29_strm0_ready         ( DownstreamStackBusLane[62][29].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane29_strm0_cntl          ( DownstreamStackBusLane[62][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane29_strm0_data          ( DownstreamStackBusLane[62][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane29_strm0_data_valid    ( DownstreamStackBusLane[62][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane29_strm1_ready         ( DownstreamStackBusLane[62][29].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane29_strm1_cntl          ( DownstreamStackBusLane[62][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane29_strm1_data          ( DownstreamStackBusLane[62][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane29_strm1_data_valid    ( DownstreamStackBusLane[62][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane30_strm0_ready         ( DownstreamStackBusLane[62][30].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane30_strm0_cntl          ( DownstreamStackBusLane[62][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane30_strm0_data          ( DownstreamStackBusLane[62][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane30_strm0_data_valid    ( DownstreamStackBusLane[62][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane30_strm1_ready         ( DownstreamStackBusLane[62][30].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane30_strm1_cntl          ( DownstreamStackBusLane[62][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane30_strm1_data          ( DownstreamStackBusLane[62][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane30_strm1_data_valid    ( DownstreamStackBusLane[62][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 62, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane31_strm0_ready         ( DownstreamStackBusLane[62][31].pe__std__lane_strm0_ready              ),      
        .std__pe62__lane31_strm0_cntl          ( DownstreamStackBusLane[62][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe62__lane31_strm0_data          ( DownstreamStackBusLane[62][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe62__lane31_strm0_data_valid    ( DownstreamStackBusLane[62][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__std__lane31_strm1_ready         ( DownstreamStackBusLane[62][31].pe__std__lane_strm1_ready              ),      
        .std__pe62__lane31_strm1_cntl          ( DownstreamStackBusLane[62][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe62__lane31_strm1_data          ( DownstreamStackBusLane[62][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe62__lane31_strm1_data_valid    ( DownstreamStackBusLane[62][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane0_strm0_ready         ( DownstreamStackBusLane[63][0].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane0_strm0_cntl          ( DownstreamStackBusLane[63][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane0_strm0_data          ( DownstreamStackBusLane[63][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane0_strm0_data_valid    ( DownstreamStackBusLane[63][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane0_strm1_ready         ( DownstreamStackBusLane[63][0].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane0_strm1_cntl          ( DownstreamStackBusLane[63][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane0_strm1_data          ( DownstreamStackBusLane[63][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane0_strm1_data_valid    ( DownstreamStackBusLane[63][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane1_strm0_ready         ( DownstreamStackBusLane[63][1].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane1_strm0_cntl          ( DownstreamStackBusLane[63][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane1_strm0_data          ( DownstreamStackBusLane[63][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane1_strm0_data_valid    ( DownstreamStackBusLane[63][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane1_strm1_ready         ( DownstreamStackBusLane[63][1].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane1_strm1_cntl          ( DownstreamStackBusLane[63][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane1_strm1_data          ( DownstreamStackBusLane[63][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane1_strm1_data_valid    ( DownstreamStackBusLane[63][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane2_strm0_ready         ( DownstreamStackBusLane[63][2].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane2_strm0_cntl          ( DownstreamStackBusLane[63][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane2_strm0_data          ( DownstreamStackBusLane[63][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane2_strm0_data_valid    ( DownstreamStackBusLane[63][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane2_strm1_ready         ( DownstreamStackBusLane[63][2].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane2_strm1_cntl          ( DownstreamStackBusLane[63][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane2_strm1_data          ( DownstreamStackBusLane[63][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane2_strm1_data_valid    ( DownstreamStackBusLane[63][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane3_strm0_ready         ( DownstreamStackBusLane[63][3].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane3_strm0_cntl          ( DownstreamStackBusLane[63][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane3_strm0_data          ( DownstreamStackBusLane[63][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane3_strm0_data_valid    ( DownstreamStackBusLane[63][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane3_strm1_ready         ( DownstreamStackBusLane[63][3].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane3_strm1_cntl          ( DownstreamStackBusLane[63][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane3_strm1_data          ( DownstreamStackBusLane[63][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane3_strm1_data_valid    ( DownstreamStackBusLane[63][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane4_strm0_ready         ( DownstreamStackBusLane[63][4].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane4_strm0_cntl          ( DownstreamStackBusLane[63][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane4_strm0_data          ( DownstreamStackBusLane[63][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane4_strm0_data_valid    ( DownstreamStackBusLane[63][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane4_strm1_ready         ( DownstreamStackBusLane[63][4].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane4_strm1_cntl          ( DownstreamStackBusLane[63][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane4_strm1_data          ( DownstreamStackBusLane[63][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane4_strm1_data_valid    ( DownstreamStackBusLane[63][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane5_strm0_ready         ( DownstreamStackBusLane[63][5].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane5_strm0_cntl          ( DownstreamStackBusLane[63][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane5_strm0_data          ( DownstreamStackBusLane[63][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane5_strm0_data_valid    ( DownstreamStackBusLane[63][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane5_strm1_ready         ( DownstreamStackBusLane[63][5].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane5_strm1_cntl          ( DownstreamStackBusLane[63][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane5_strm1_data          ( DownstreamStackBusLane[63][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane5_strm1_data_valid    ( DownstreamStackBusLane[63][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane6_strm0_ready         ( DownstreamStackBusLane[63][6].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane6_strm0_cntl          ( DownstreamStackBusLane[63][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane6_strm0_data          ( DownstreamStackBusLane[63][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane6_strm0_data_valid    ( DownstreamStackBusLane[63][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane6_strm1_ready         ( DownstreamStackBusLane[63][6].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane6_strm1_cntl          ( DownstreamStackBusLane[63][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane6_strm1_data          ( DownstreamStackBusLane[63][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane6_strm1_data_valid    ( DownstreamStackBusLane[63][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane7_strm0_ready         ( DownstreamStackBusLane[63][7].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane7_strm0_cntl          ( DownstreamStackBusLane[63][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane7_strm0_data          ( DownstreamStackBusLane[63][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane7_strm0_data_valid    ( DownstreamStackBusLane[63][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane7_strm1_ready         ( DownstreamStackBusLane[63][7].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane7_strm1_cntl          ( DownstreamStackBusLane[63][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane7_strm1_data          ( DownstreamStackBusLane[63][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane7_strm1_data_valid    ( DownstreamStackBusLane[63][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane8_strm0_ready         ( DownstreamStackBusLane[63][8].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane8_strm0_cntl          ( DownstreamStackBusLane[63][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane8_strm0_data          ( DownstreamStackBusLane[63][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane8_strm0_data_valid    ( DownstreamStackBusLane[63][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane8_strm1_ready         ( DownstreamStackBusLane[63][8].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane8_strm1_cntl          ( DownstreamStackBusLane[63][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane8_strm1_data          ( DownstreamStackBusLane[63][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane8_strm1_data_valid    ( DownstreamStackBusLane[63][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane9_strm0_ready         ( DownstreamStackBusLane[63][9].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane9_strm0_cntl          ( DownstreamStackBusLane[63][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane9_strm0_data          ( DownstreamStackBusLane[63][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane9_strm0_data_valid    ( DownstreamStackBusLane[63][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane9_strm1_ready         ( DownstreamStackBusLane[63][9].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane9_strm1_cntl          ( DownstreamStackBusLane[63][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane9_strm1_data          ( DownstreamStackBusLane[63][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane9_strm1_data_valid    ( DownstreamStackBusLane[63][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane10_strm0_ready         ( DownstreamStackBusLane[63][10].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane10_strm0_cntl          ( DownstreamStackBusLane[63][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane10_strm0_data          ( DownstreamStackBusLane[63][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane10_strm0_data_valid    ( DownstreamStackBusLane[63][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane10_strm1_ready         ( DownstreamStackBusLane[63][10].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane10_strm1_cntl          ( DownstreamStackBusLane[63][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane10_strm1_data          ( DownstreamStackBusLane[63][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane10_strm1_data_valid    ( DownstreamStackBusLane[63][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane11_strm0_ready         ( DownstreamStackBusLane[63][11].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane11_strm0_cntl          ( DownstreamStackBusLane[63][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane11_strm0_data          ( DownstreamStackBusLane[63][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane11_strm0_data_valid    ( DownstreamStackBusLane[63][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane11_strm1_ready         ( DownstreamStackBusLane[63][11].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane11_strm1_cntl          ( DownstreamStackBusLane[63][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane11_strm1_data          ( DownstreamStackBusLane[63][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane11_strm1_data_valid    ( DownstreamStackBusLane[63][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane12_strm0_ready         ( DownstreamStackBusLane[63][12].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane12_strm0_cntl          ( DownstreamStackBusLane[63][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane12_strm0_data          ( DownstreamStackBusLane[63][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane12_strm0_data_valid    ( DownstreamStackBusLane[63][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane12_strm1_ready         ( DownstreamStackBusLane[63][12].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane12_strm1_cntl          ( DownstreamStackBusLane[63][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane12_strm1_data          ( DownstreamStackBusLane[63][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane12_strm1_data_valid    ( DownstreamStackBusLane[63][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane13_strm0_ready         ( DownstreamStackBusLane[63][13].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane13_strm0_cntl          ( DownstreamStackBusLane[63][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane13_strm0_data          ( DownstreamStackBusLane[63][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane13_strm0_data_valid    ( DownstreamStackBusLane[63][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane13_strm1_ready         ( DownstreamStackBusLane[63][13].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane13_strm1_cntl          ( DownstreamStackBusLane[63][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane13_strm1_data          ( DownstreamStackBusLane[63][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane13_strm1_data_valid    ( DownstreamStackBusLane[63][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane14_strm0_ready         ( DownstreamStackBusLane[63][14].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane14_strm0_cntl          ( DownstreamStackBusLane[63][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane14_strm0_data          ( DownstreamStackBusLane[63][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane14_strm0_data_valid    ( DownstreamStackBusLane[63][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane14_strm1_ready         ( DownstreamStackBusLane[63][14].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane14_strm1_cntl          ( DownstreamStackBusLane[63][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane14_strm1_data          ( DownstreamStackBusLane[63][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane14_strm1_data_valid    ( DownstreamStackBusLane[63][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane15_strm0_ready         ( DownstreamStackBusLane[63][15].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane15_strm0_cntl          ( DownstreamStackBusLane[63][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane15_strm0_data          ( DownstreamStackBusLane[63][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane15_strm0_data_valid    ( DownstreamStackBusLane[63][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane15_strm1_ready         ( DownstreamStackBusLane[63][15].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane15_strm1_cntl          ( DownstreamStackBusLane[63][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane15_strm1_data          ( DownstreamStackBusLane[63][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane15_strm1_data_valid    ( DownstreamStackBusLane[63][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane16_strm0_ready         ( DownstreamStackBusLane[63][16].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane16_strm0_cntl          ( DownstreamStackBusLane[63][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane16_strm0_data          ( DownstreamStackBusLane[63][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane16_strm0_data_valid    ( DownstreamStackBusLane[63][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane16_strm1_ready         ( DownstreamStackBusLane[63][16].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane16_strm1_cntl          ( DownstreamStackBusLane[63][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane16_strm1_data          ( DownstreamStackBusLane[63][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane16_strm1_data_valid    ( DownstreamStackBusLane[63][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane17_strm0_ready         ( DownstreamStackBusLane[63][17].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane17_strm0_cntl          ( DownstreamStackBusLane[63][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane17_strm0_data          ( DownstreamStackBusLane[63][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane17_strm0_data_valid    ( DownstreamStackBusLane[63][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane17_strm1_ready         ( DownstreamStackBusLane[63][17].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane17_strm1_cntl          ( DownstreamStackBusLane[63][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane17_strm1_data          ( DownstreamStackBusLane[63][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane17_strm1_data_valid    ( DownstreamStackBusLane[63][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane18_strm0_ready         ( DownstreamStackBusLane[63][18].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane18_strm0_cntl          ( DownstreamStackBusLane[63][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane18_strm0_data          ( DownstreamStackBusLane[63][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane18_strm0_data_valid    ( DownstreamStackBusLane[63][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane18_strm1_ready         ( DownstreamStackBusLane[63][18].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane18_strm1_cntl          ( DownstreamStackBusLane[63][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane18_strm1_data          ( DownstreamStackBusLane[63][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane18_strm1_data_valid    ( DownstreamStackBusLane[63][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane19_strm0_ready         ( DownstreamStackBusLane[63][19].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane19_strm0_cntl          ( DownstreamStackBusLane[63][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane19_strm0_data          ( DownstreamStackBusLane[63][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane19_strm0_data_valid    ( DownstreamStackBusLane[63][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane19_strm1_ready         ( DownstreamStackBusLane[63][19].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane19_strm1_cntl          ( DownstreamStackBusLane[63][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane19_strm1_data          ( DownstreamStackBusLane[63][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane19_strm1_data_valid    ( DownstreamStackBusLane[63][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane20_strm0_ready         ( DownstreamStackBusLane[63][20].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane20_strm0_cntl          ( DownstreamStackBusLane[63][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane20_strm0_data          ( DownstreamStackBusLane[63][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane20_strm0_data_valid    ( DownstreamStackBusLane[63][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane20_strm1_ready         ( DownstreamStackBusLane[63][20].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane20_strm1_cntl          ( DownstreamStackBusLane[63][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane20_strm1_data          ( DownstreamStackBusLane[63][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane20_strm1_data_valid    ( DownstreamStackBusLane[63][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane21_strm0_ready         ( DownstreamStackBusLane[63][21].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane21_strm0_cntl          ( DownstreamStackBusLane[63][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane21_strm0_data          ( DownstreamStackBusLane[63][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane21_strm0_data_valid    ( DownstreamStackBusLane[63][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane21_strm1_ready         ( DownstreamStackBusLane[63][21].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane21_strm1_cntl          ( DownstreamStackBusLane[63][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane21_strm1_data          ( DownstreamStackBusLane[63][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane21_strm1_data_valid    ( DownstreamStackBusLane[63][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane22_strm0_ready         ( DownstreamStackBusLane[63][22].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane22_strm0_cntl          ( DownstreamStackBusLane[63][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane22_strm0_data          ( DownstreamStackBusLane[63][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane22_strm0_data_valid    ( DownstreamStackBusLane[63][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane22_strm1_ready         ( DownstreamStackBusLane[63][22].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane22_strm1_cntl          ( DownstreamStackBusLane[63][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane22_strm1_data          ( DownstreamStackBusLane[63][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane22_strm1_data_valid    ( DownstreamStackBusLane[63][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane23_strm0_ready         ( DownstreamStackBusLane[63][23].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane23_strm0_cntl          ( DownstreamStackBusLane[63][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane23_strm0_data          ( DownstreamStackBusLane[63][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane23_strm0_data_valid    ( DownstreamStackBusLane[63][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane23_strm1_ready         ( DownstreamStackBusLane[63][23].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane23_strm1_cntl          ( DownstreamStackBusLane[63][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane23_strm1_data          ( DownstreamStackBusLane[63][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane23_strm1_data_valid    ( DownstreamStackBusLane[63][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane24_strm0_ready         ( DownstreamStackBusLane[63][24].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane24_strm0_cntl          ( DownstreamStackBusLane[63][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane24_strm0_data          ( DownstreamStackBusLane[63][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane24_strm0_data_valid    ( DownstreamStackBusLane[63][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane24_strm1_ready         ( DownstreamStackBusLane[63][24].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane24_strm1_cntl          ( DownstreamStackBusLane[63][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane24_strm1_data          ( DownstreamStackBusLane[63][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane24_strm1_data_valid    ( DownstreamStackBusLane[63][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane25_strm0_ready         ( DownstreamStackBusLane[63][25].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane25_strm0_cntl          ( DownstreamStackBusLane[63][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane25_strm0_data          ( DownstreamStackBusLane[63][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane25_strm0_data_valid    ( DownstreamStackBusLane[63][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane25_strm1_ready         ( DownstreamStackBusLane[63][25].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane25_strm1_cntl          ( DownstreamStackBusLane[63][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane25_strm1_data          ( DownstreamStackBusLane[63][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane25_strm1_data_valid    ( DownstreamStackBusLane[63][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane26_strm0_ready         ( DownstreamStackBusLane[63][26].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane26_strm0_cntl          ( DownstreamStackBusLane[63][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane26_strm0_data          ( DownstreamStackBusLane[63][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane26_strm0_data_valid    ( DownstreamStackBusLane[63][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane26_strm1_ready         ( DownstreamStackBusLane[63][26].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane26_strm1_cntl          ( DownstreamStackBusLane[63][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane26_strm1_data          ( DownstreamStackBusLane[63][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane26_strm1_data_valid    ( DownstreamStackBusLane[63][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane27_strm0_ready         ( DownstreamStackBusLane[63][27].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane27_strm0_cntl          ( DownstreamStackBusLane[63][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane27_strm0_data          ( DownstreamStackBusLane[63][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane27_strm0_data_valid    ( DownstreamStackBusLane[63][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane27_strm1_ready         ( DownstreamStackBusLane[63][27].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane27_strm1_cntl          ( DownstreamStackBusLane[63][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane27_strm1_data          ( DownstreamStackBusLane[63][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane27_strm1_data_valid    ( DownstreamStackBusLane[63][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane28_strm0_ready         ( DownstreamStackBusLane[63][28].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane28_strm0_cntl          ( DownstreamStackBusLane[63][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane28_strm0_data          ( DownstreamStackBusLane[63][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane28_strm0_data_valid    ( DownstreamStackBusLane[63][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane28_strm1_ready         ( DownstreamStackBusLane[63][28].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane28_strm1_cntl          ( DownstreamStackBusLane[63][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane28_strm1_data          ( DownstreamStackBusLane[63][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane28_strm1_data_valid    ( DownstreamStackBusLane[63][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane29_strm0_ready         ( DownstreamStackBusLane[63][29].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane29_strm0_cntl          ( DownstreamStackBusLane[63][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane29_strm0_data          ( DownstreamStackBusLane[63][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane29_strm0_data_valid    ( DownstreamStackBusLane[63][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane29_strm1_ready         ( DownstreamStackBusLane[63][29].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane29_strm1_cntl          ( DownstreamStackBusLane[63][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane29_strm1_data          ( DownstreamStackBusLane[63][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane29_strm1_data_valid    ( DownstreamStackBusLane[63][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane30_strm0_ready         ( DownstreamStackBusLane[63][30].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane30_strm0_cntl          ( DownstreamStackBusLane[63][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane30_strm0_data          ( DownstreamStackBusLane[63][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane30_strm0_data_valid    ( DownstreamStackBusLane[63][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane30_strm1_ready         ( DownstreamStackBusLane[63][30].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane30_strm1_cntl          ( DownstreamStackBusLane[63][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane30_strm1_data          ( DownstreamStackBusLane[63][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane30_strm1_data_valid    ( DownstreamStackBusLane[63][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 63, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane31_strm0_ready         ( DownstreamStackBusLane[63][31].pe__std__lane_strm0_ready              ),      
        .std__pe63__lane31_strm0_cntl          ( DownstreamStackBusLane[63][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe63__lane31_strm0_data          ( DownstreamStackBusLane[63][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe63__lane31_strm0_data_valid    ( DownstreamStackBusLane[63][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__std__lane31_strm1_ready         ( DownstreamStackBusLane[63][31].pe__std__lane_strm1_ready              ),      
        .std__pe63__lane31_strm1_cntl          ( DownstreamStackBusLane[63][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe63__lane31_strm1_data          ( DownstreamStackBusLane[63][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe63__lane31_strm1_data_valid    ( DownstreamStackBusLane[63][31].cb_test.std__pe__lane_strm1_data_valid ),      
        