
  // lane0 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane0_toStOp_strm_cntl                 ;
  reg                                                         lane0_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane0_toStOp_strm_data                 ;
  reg                                                         lane0_toStOp_strm_fifo_write           ;
  wire                                                        lane0_toStOp_strm_ready                ;
  wire                                                        lane0_toStOp_strm_fifo_read            ;
  reg                                                         lane0_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane0_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane0_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane0_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane0_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane0_toStOp_strm_fifo_read_data       ;
  wire                                                        lane0_toStOp_strm_fifo_data_available  ;
  // lane1 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane1_toStOp_strm_cntl                 ;
  reg                                                         lane1_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane1_toStOp_strm_data                 ;
  reg                                                         lane1_toStOp_strm_fifo_write           ;
  wire                                                        lane1_toStOp_strm_ready                ;
  wire                                                        lane1_toStOp_strm_fifo_read            ;
  reg                                                         lane1_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane1_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane1_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane1_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane1_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane1_toStOp_strm_fifo_read_data       ;
  wire                                                        lane1_toStOp_strm_fifo_data_available  ;
  // lane2 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane2_toStOp_strm_cntl                 ;
  reg                                                         lane2_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane2_toStOp_strm_data                 ;
  reg                                                         lane2_toStOp_strm_fifo_write           ;
  wire                                                        lane2_toStOp_strm_ready                ;
  wire                                                        lane2_toStOp_strm_fifo_read            ;
  reg                                                         lane2_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane2_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane2_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane2_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane2_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane2_toStOp_strm_fifo_read_data       ;
  wire                                                        lane2_toStOp_strm_fifo_data_available  ;
  // lane3 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane3_toStOp_strm_cntl                 ;
  reg                                                         lane3_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane3_toStOp_strm_data                 ;
  reg                                                         lane3_toStOp_strm_fifo_write           ;
  wire                                                        lane3_toStOp_strm_ready                ;
  wire                                                        lane3_toStOp_strm_fifo_read            ;
  reg                                                         lane3_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane3_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane3_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane3_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane3_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane3_toStOp_strm_fifo_read_data       ;
  wire                                                        lane3_toStOp_strm_fifo_data_available  ;
  // lane4 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane4_toStOp_strm_cntl                 ;
  reg                                                         lane4_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane4_toStOp_strm_data                 ;
  reg                                                         lane4_toStOp_strm_fifo_write           ;
  wire                                                        lane4_toStOp_strm_ready                ;
  wire                                                        lane4_toStOp_strm_fifo_read            ;
  reg                                                         lane4_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane4_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane4_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane4_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane4_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane4_toStOp_strm_fifo_read_data       ;
  wire                                                        lane4_toStOp_strm_fifo_data_available  ;
  // lane5 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane5_toStOp_strm_cntl                 ;
  reg                                                         lane5_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane5_toStOp_strm_data                 ;
  reg                                                         lane5_toStOp_strm_fifo_write           ;
  wire                                                        lane5_toStOp_strm_ready                ;
  wire                                                        lane5_toStOp_strm_fifo_read            ;
  reg                                                         lane5_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane5_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane5_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane5_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane5_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane5_toStOp_strm_fifo_read_data       ;
  wire                                                        lane5_toStOp_strm_fifo_data_available  ;
  // lane6 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane6_toStOp_strm_cntl                 ;
  reg                                                         lane6_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane6_toStOp_strm_data                 ;
  reg                                                         lane6_toStOp_strm_fifo_write           ;
  wire                                                        lane6_toStOp_strm_ready                ;
  wire                                                        lane6_toStOp_strm_fifo_read            ;
  reg                                                         lane6_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane6_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane6_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane6_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane6_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane6_toStOp_strm_fifo_read_data       ;
  wire                                                        lane6_toStOp_strm_fifo_data_available  ;
  // lane7 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane7_toStOp_strm_cntl                 ;
  reg                                                         lane7_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane7_toStOp_strm_data                 ;
  reg                                                         lane7_toStOp_strm_fifo_write           ;
  wire                                                        lane7_toStOp_strm_ready                ;
  wire                                                        lane7_toStOp_strm_fifo_read            ;
  reg                                                         lane7_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane7_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane7_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane7_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane7_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane7_toStOp_strm_fifo_read_data       ;
  wire                                                        lane7_toStOp_strm_fifo_data_available  ;
  // lane8 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane8_toStOp_strm_cntl                 ;
  reg                                                         lane8_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane8_toStOp_strm_data                 ;
  reg                                                         lane8_toStOp_strm_fifo_write           ;
  wire                                                        lane8_toStOp_strm_ready                ;
  wire                                                        lane8_toStOp_strm_fifo_read            ;
  reg                                                         lane8_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane8_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane8_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane8_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane8_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane8_toStOp_strm_fifo_read_data       ;
  wire                                                        lane8_toStOp_strm_fifo_data_available  ;
  // lane9 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane9_toStOp_strm_cntl                 ;
  reg                                                         lane9_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane9_toStOp_strm_data                 ;
  reg                                                         lane9_toStOp_strm_fifo_write           ;
  wire                                                        lane9_toStOp_strm_ready                ;
  wire                                                        lane9_toStOp_strm_fifo_read            ;
  reg                                                         lane9_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane9_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane9_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane9_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane9_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane9_toStOp_strm_fifo_read_data       ;
  wire                                                        lane9_toStOp_strm_fifo_data_available  ;
  // lane10 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane10_toStOp_strm_cntl                 ;
  reg                                                         lane10_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane10_toStOp_strm_data                 ;
  reg                                                         lane10_toStOp_strm_fifo_write           ;
  wire                                                        lane10_toStOp_strm_ready                ;
  wire                                                        lane10_toStOp_strm_fifo_read            ;
  reg                                                         lane10_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane10_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane10_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane10_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane10_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane10_toStOp_strm_fifo_read_data       ;
  wire                                                        lane10_toStOp_strm_fifo_data_available  ;
  // lane11 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane11_toStOp_strm_cntl                 ;
  reg                                                         lane11_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane11_toStOp_strm_data                 ;
  reg                                                         lane11_toStOp_strm_fifo_write           ;
  wire                                                        lane11_toStOp_strm_ready                ;
  wire                                                        lane11_toStOp_strm_fifo_read            ;
  reg                                                         lane11_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane11_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane11_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane11_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane11_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane11_toStOp_strm_fifo_read_data       ;
  wire                                                        lane11_toStOp_strm_fifo_data_available  ;
  // lane12 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane12_toStOp_strm_cntl                 ;
  reg                                                         lane12_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane12_toStOp_strm_data                 ;
  reg                                                         lane12_toStOp_strm_fifo_write           ;
  wire                                                        lane12_toStOp_strm_ready                ;
  wire                                                        lane12_toStOp_strm_fifo_read            ;
  reg                                                         lane12_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane12_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane12_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane12_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane12_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane12_toStOp_strm_fifo_read_data       ;
  wire                                                        lane12_toStOp_strm_fifo_data_available  ;
  // lane13 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane13_toStOp_strm_cntl                 ;
  reg                                                         lane13_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane13_toStOp_strm_data                 ;
  reg                                                         lane13_toStOp_strm_fifo_write           ;
  wire                                                        lane13_toStOp_strm_ready                ;
  wire                                                        lane13_toStOp_strm_fifo_read            ;
  reg                                                         lane13_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane13_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane13_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane13_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane13_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane13_toStOp_strm_fifo_read_data       ;
  wire                                                        lane13_toStOp_strm_fifo_data_available  ;
  // lane14 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane14_toStOp_strm_cntl                 ;
  reg                                                         lane14_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane14_toStOp_strm_data                 ;
  reg                                                         lane14_toStOp_strm_fifo_write           ;
  wire                                                        lane14_toStOp_strm_ready                ;
  wire                                                        lane14_toStOp_strm_fifo_read            ;
  reg                                                         lane14_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane14_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane14_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane14_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane14_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane14_toStOp_strm_fifo_read_data       ;
  wire                                                        lane14_toStOp_strm_fifo_data_available  ;
  // lane15 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane15_toStOp_strm_cntl                 ;
  reg                                                         lane15_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane15_toStOp_strm_data                 ;
  reg                                                         lane15_toStOp_strm_fifo_write           ;
  wire                                                        lane15_toStOp_strm_ready                ;
  wire                                                        lane15_toStOp_strm_fifo_read            ;
  reg                                                         lane15_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane15_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane15_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane15_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane15_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane15_toStOp_strm_fifo_read_data       ;
  wire                                                        lane15_toStOp_strm_fifo_data_available  ;
  // lane16 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane16_toStOp_strm_cntl                 ;
  reg                                                         lane16_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane16_toStOp_strm_data                 ;
  reg                                                         lane16_toStOp_strm_fifo_write           ;
  wire                                                        lane16_toStOp_strm_ready                ;
  wire                                                        lane16_toStOp_strm_fifo_read            ;
  reg                                                         lane16_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane16_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane16_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane16_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane16_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane16_toStOp_strm_fifo_read_data       ;
  wire                                                        lane16_toStOp_strm_fifo_data_available  ;
  // lane17 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane17_toStOp_strm_cntl                 ;
  reg                                                         lane17_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane17_toStOp_strm_data                 ;
  reg                                                         lane17_toStOp_strm_fifo_write           ;
  wire                                                        lane17_toStOp_strm_ready                ;
  wire                                                        lane17_toStOp_strm_fifo_read            ;
  reg                                                         lane17_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane17_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane17_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane17_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane17_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane17_toStOp_strm_fifo_read_data       ;
  wire                                                        lane17_toStOp_strm_fifo_data_available  ;
  // lane18 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane18_toStOp_strm_cntl                 ;
  reg                                                         lane18_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane18_toStOp_strm_data                 ;
  reg                                                         lane18_toStOp_strm_fifo_write           ;
  wire                                                        lane18_toStOp_strm_ready                ;
  wire                                                        lane18_toStOp_strm_fifo_read            ;
  reg                                                         lane18_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane18_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane18_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane18_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane18_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane18_toStOp_strm_fifo_read_data       ;
  wire                                                        lane18_toStOp_strm_fifo_data_available  ;
  // lane19 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane19_toStOp_strm_cntl                 ;
  reg                                                         lane19_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane19_toStOp_strm_data                 ;
  reg                                                         lane19_toStOp_strm_fifo_write           ;
  wire                                                        lane19_toStOp_strm_ready                ;
  wire                                                        lane19_toStOp_strm_fifo_read            ;
  reg                                                         lane19_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane19_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane19_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane19_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane19_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane19_toStOp_strm_fifo_read_data       ;
  wire                                                        lane19_toStOp_strm_fifo_data_available  ;
  // lane20 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane20_toStOp_strm_cntl                 ;
  reg                                                         lane20_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane20_toStOp_strm_data                 ;
  reg                                                         lane20_toStOp_strm_fifo_write           ;
  wire                                                        lane20_toStOp_strm_ready                ;
  wire                                                        lane20_toStOp_strm_fifo_read            ;
  reg                                                         lane20_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane20_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane20_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane20_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane20_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane20_toStOp_strm_fifo_read_data       ;
  wire                                                        lane20_toStOp_strm_fifo_data_available  ;
  // lane21 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane21_toStOp_strm_cntl                 ;
  reg                                                         lane21_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane21_toStOp_strm_data                 ;
  reg                                                         lane21_toStOp_strm_fifo_write           ;
  wire                                                        lane21_toStOp_strm_ready                ;
  wire                                                        lane21_toStOp_strm_fifo_read            ;
  reg                                                         lane21_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane21_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane21_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane21_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane21_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane21_toStOp_strm_fifo_read_data       ;
  wire                                                        lane21_toStOp_strm_fifo_data_available  ;
  // lane22 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane22_toStOp_strm_cntl                 ;
  reg                                                         lane22_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane22_toStOp_strm_data                 ;
  reg                                                         lane22_toStOp_strm_fifo_write           ;
  wire                                                        lane22_toStOp_strm_ready                ;
  wire                                                        lane22_toStOp_strm_fifo_read            ;
  reg                                                         lane22_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane22_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane22_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane22_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane22_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane22_toStOp_strm_fifo_read_data       ;
  wire                                                        lane22_toStOp_strm_fifo_data_available  ;
  // lane23 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane23_toStOp_strm_cntl                 ;
  reg                                                         lane23_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane23_toStOp_strm_data                 ;
  reg                                                         lane23_toStOp_strm_fifo_write           ;
  wire                                                        lane23_toStOp_strm_ready                ;
  wire                                                        lane23_toStOp_strm_fifo_read            ;
  reg                                                         lane23_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane23_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane23_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane23_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane23_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane23_toStOp_strm_fifo_read_data       ;
  wire                                                        lane23_toStOp_strm_fifo_data_available  ;
  // lane24 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane24_toStOp_strm_cntl                 ;
  reg                                                         lane24_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane24_toStOp_strm_data                 ;
  reg                                                         lane24_toStOp_strm_fifo_write           ;
  wire                                                        lane24_toStOp_strm_ready                ;
  wire                                                        lane24_toStOp_strm_fifo_read            ;
  reg                                                         lane24_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane24_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane24_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane24_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane24_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane24_toStOp_strm_fifo_read_data       ;
  wire                                                        lane24_toStOp_strm_fifo_data_available  ;
  // lane25 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane25_toStOp_strm_cntl                 ;
  reg                                                         lane25_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane25_toStOp_strm_data                 ;
  reg                                                         lane25_toStOp_strm_fifo_write           ;
  wire                                                        lane25_toStOp_strm_ready                ;
  wire                                                        lane25_toStOp_strm_fifo_read            ;
  reg                                                         lane25_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane25_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane25_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane25_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane25_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane25_toStOp_strm_fifo_read_data       ;
  wire                                                        lane25_toStOp_strm_fifo_data_available  ;
  // lane26 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane26_toStOp_strm_cntl                 ;
  reg                                                         lane26_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane26_toStOp_strm_data                 ;
  reg                                                         lane26_toStOp_strm_fifo_write           ;
  wire                                                        lane26_toStOp_strm_ready                ;
  wire                                                        lane26_toStOp_strm_fifo_read            ;
  reg                                                         lane26_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane26_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane26_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane26_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane26_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane26_toStOp_strm_fifo_read_data       ;
  wire                                                        lane26_toStOp_strm_fifo_data_available  ;
  // lane27 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane27_toStOp_strm_cntl                 ;
  reg                                                         lane27_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane27_toStOp_strm_data                 ;
  reg                                                         lane27_toStOp_strm_fifo_write           ;
  wire                                                        lane27_toStOp_strm_ready                ;
  wire                                                        lane27_toStOp_strm_fifo_read            ;
  reg                                                         lane27_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane27_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane27_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane27_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane27_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane27_toStOp_strm_fifo_read_data       ;
  wire                                                        lane27_toStOp_strm_fifo_data_available  ;
  // lane28 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane28_toStOp_strm_cntl                 ;
  reg                                                         lane28_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane28_toStOp_strm_data                 ;
  reg                                                         lane28_toStOp_strm_fifo_write           ;
  wire                                                        lane28_toStOp_strm_ready                ;
  wire                                                        lane28_toStOp_strm_fifo_read            ;
  reg                                                         lane28_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane28_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane28_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane28_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane28_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane28_toStOp_strm_fifo_read_data       ;
  wire                                                        lane28_toStOp_strm_fifo_data_available  ;
  // lane29 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane29_toStOp_strm_cntl                 ;
  reg                                                         lane29_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane29_toStOp_strm_data                 ;
  reg                                                         lane29_toStOp_strm_fifo_write           ;
  wire                                                        lane29_toStOp_strm_ready                ;
  wire                                                        lane29_toStOp_strm_fifo_read            ;
  reg                                                         lane29_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane29_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane29_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane29_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane29_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane29_toStOp_strm_fifo_read_data       ;
  wire                                                        lane29_toStOp_strm_fifo_data_available  ;
  // lane30 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane30_toStOp_strm_cntl                 ;
  reg                                                         lane30_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane30_toStOp_strm_data                 ;
  reg                                                         lane30_toStOp_strm_fifo_write           ;
  wire                                                        lane30_toStOp_strm_ready                ;
  wire                                                        lane30_toStOp_strm_fifo_read            ;
  reg                                                         lane30_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane30_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane30_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane30_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane30_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane30_toStOp_strm_fifo_read_data       ;
  wire                                                        lane30_toStOp_strm_fifo_data_available  ;
  // lane31 to NoC 
  reg  [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane31_toStOp_strm_cntl                 ;
  reg                                                         lane31_toStOp_strm_id                   ;
  reg  [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane31_toStOp_strm_data                 ;
  reg                                                         lane31_toStOp_strm_fifo_write           ;
  wire                                                        lane31_toStOp_strm_ready                ;
  wire                                                        lane31_toStOp_strm_fifo_read            ;
  reg                                                         lane31_toStOp_strm_fifo_read_valid      ;
  wire                                                        lane31_toStOp_strm_fifo_empty           ;
  wire [`STREAMING_OP_CNTL_STOP_TO_NOC_FIFO_EOP_COUNT_RANGE ] lane31_toStOp_strm_fifo_eop_count       ;
  wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE                  ] lane31_toStOp_strm_fifo_read_cntl       ;
  wire                                                        lane31_toStOp_strm_fifo_read_id         ;
  wire [`STREAMING_OP_CNTL_DATA_RANGE                       ] lane31_toStOp_strm_fifo_read_data       ;
  wire                                                        lane31_toStOp_strm_fifo_data_available  ;