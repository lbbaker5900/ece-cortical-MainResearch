
               // OOB carries PE configuration                                               
               .sti__cntl__oob_cntl                  ( sti__cntl__oob_cntl               ),      
               .sti__cntl__oob_valid                 ( sti__cntl__oob_valid              ),      
               .cntl__sti__oob_ready                 ( cntl__sti__oob_ready              ),      
               .sti__cntl__oob_type                  ( sti__cntl__oob_type               ),      
               .sti__cntl__oob_data                  ( sti__cntl__oob_data               ),      