
  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe0__allSynchronized    ( GenStackBus[0].sys__pe__allSynchronized           ), 
        .pe0__sys__thisSynchronized   ( GenStackBus[0].pe__sys__thisSynchronized          ), 
        .pe0__sys__ready              ( GenStackBus[0].pe__sys__ready                     ), 
        .pe0__sys__complete           ( GenStackBus[0].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe1__allSynchronized    ( GenStackBus[1].sys__pe__allSynchronized           ), 
        .pe1__sys__thisSynchronized   ( GenStackBus[1].pe__sys__thisSynchronized          ), 
        .pe1__sys__ready              ( GenStackBus[1].pe__sys__ready                     ), 
        .pe1__sys__complete           ( GenStackBus[1].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe2__allSynchronized    ( GenStackBus[2].sys__pe__allSynchronized           ), 
        .pe2__sys__thisSynchronized   ( GenStackBus[2].pe__sys__thisSynchronized          ), 
        .pe2__sys__ready              ( GenStackBus[2].pe__sys__ready                     ), 
        .pe2__sys__complete           ( GenStackBus[2].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe3__allSynchronized    ( GenStackBus[3].sys__pe__allSynchronized           ), 
        .pe3__sys__thisSynchronized   ( GenStackBus[3].pe__sys__thisSynchronized          ), 
        .pe3__sys__ready              ( GenStackBus[3].pe__sys__ready                     ), 
        .pe3__sys__complete           ( GenStackBus[3].pe__sys__complete                  ), 
