
    assign reg__scntl__lane0_ready = reg__scntl__ready [0]    ;
    assign scntl__reg__valid [0]   = scntl__reg__lane0_valid  ;
    assign scntl__reg__data  [0]   = scntl__reg__lane0_data   ;

    assign reg__scntl__lane1_ready = reg__scntl__ready [1]    ;
    assign scntl__reg__valid [1]   = scntl__reg__lane1_valid  ;
    assign scntl__reg__data  [1]   = scntl__reg__lane1_data   ;

    assign reg__scntl__lane2_ready = reg__scntl__ready [2]    ;
    assign scntl__reg__valid [2]   = scntl__reg__lane2_valid  ;
    assign scntl__reg__data  [2]   = scntl__reg__lane2_data   ;

    assign reg__scntl__lane3_ready = reg__scntl__ready [3]    ;
    assign scntl__reg__valid [3]   = scntl__reg__lane3_valid  ;
    assign scntl__reg__data  [3]   = scntl__reg__lane3_data   ;

    assign reg__scntl__lane4_ready = reg__scntl__ready [4]    ;
    assign scntl__reg__valid [4]   = scntl__reg__lane4_valid  ;
    assign scntl__reg__data  [4]   = scntl__reg__lane4_data   ;

    assign reg__scntl__lane5_ready = reg__scntl__ready [5]    ;
    assign scntl__reg__valid [5]   = scntl__reg__lane5_valid  ;
    assign scntl__reg__data  [5]   = scntl__reg__lane5_data   ;

    assign reg__scntl__lane6_ready = reg__scntl__ready [6]    ;
    assign scntl__reg__valid [6]   = scntl__reg__lane6_valid  ;
    assign scntl__reg__data  [6]   = scntl__reg__lane6_data   ;

    assign reg__scntl__lane7_ready = reg__scntl__ready [7]    ;
    assign scntl__reg__valid [7]   = scntl__reg__lane7_valid  ;
    assign scntl__reg__data  [7]   = scntl__reg__lane7_data   ;

    assign reg__scntl__lane8_ready = reg__scntl__ready [8]    ;
    assign scntl__reg__valid [8]   = scntl__reg__lane8_valid  ;
    assign scntl__reg__data  [8]   = scntl__reg__lane8_data   ;

    assign reg__scntl__lane9_ready = reg__scntl__ready [9]    ;
    assign scntl__reg__valid [9]   = scntl__reg__lane9_valid  ;
    assign scntl__reg__data  [9]   = scntl__reg__lane9_data   ;

    assign reg__scntl__lane10_ready = reg__scntl__ready [10]    ;
    assign scntl__reg__valid [10]   = scntl__reg__lane10_valid  ;
    assign scntl__reg__data  [10]   = scntl__reg__lane10_data   ;

    assign reg__scntl__lane11_ready = reg__scntl__ready [11]    ;
    assign scntl__reg__valid [11]   = scntl__reg__lane11_valid  ;
    assign scntl__reg__data  [11]   = scntl__reg__lane11_data   ;

    assign reg__scntl__lane12_ready = reg__scntl__ready [12]    ;
    assign scntl__reg__valid [12]   = scntl__reg__lane12_valid  ;
    assign scntl__reg__data  [12]   = scntl__reg__lane12_data   ;

    assign reg__scntl__lane13_ready = reg__scntl__ready [13]    ;
    assign scntl__reg__valid [13]   = scntl__reg__lane13_valid  ;
    assign scntl__reg__data  [13]   = scntl__reg__lane13_data   ;

    assign reg__scntl__lane14_ready = reg__scntl__ready [14]    ;
    assign scntl__reg__valid [14]   = scntl__reg__lane14_valid  ;
    assign scntl__reg__data  [14]   = scntl__reg__lane14_data   ;

    assign reg__scntl__lane15_ready = reg__scntl__ready [15]    ;
    assign scntl__reg__valid [15]   = scntl__reg__lane15_valid  ;
    assign scntl__reg__data  [15]   = scntl__reg__lane15_data   ;

    assign reg__scntl__lane16_ready = reg__scntl__ready [16]    ;
    assign scntl__reg__valid [16]   = scntl__reg__lane16_valid  ;
    assign scntl__reg__data  [16]   = scntl__reg__lane16_data   ;

    assign reg__scntl__lane17_ready = reg__scntl__ready [17]    ;
    assign scntl__reg__valid [17]   = scntl__reg__lane17_valid  ;
    assign scntl__reg__data  [17]   = scntl__reg__lane17_data   ;

    assign reg__scntl__lane18_ready = reg__scntl__ready [18]    ;
    assign scntl__reg__valid [18]   = scntl__reg__lane18_valid  ;
    assign scntl__reg__data  [18]   = scntl__reg__lane18_data   ;

    assign reg__scntl__lane19_ready = reg__scntl__ready [19]    ;
    assign scntl__reg__valid [19]   = scntl__reg__lane19_valid  ;
    assign scntl__reg__data  [19]   = scntl__reg__lane19_data   ;

    assign reg__scntl__lane20_ready = reg__scntl__ready [20]    ;
    assign scntl__reg__valid [20]   = scntl__reg__lane20_valid  ;
    assign scntl__reg__data  [20]   = scntl__reg__lane20_data   ;

    assign reg__scntl__lane21_ready = reg__scntl__ready [21]    ;
    assign scntl__reg__valid [21]   = scntl__reg__lane21_valid  ;
    assign scntl__reg__data  [21]   = scntl__reg__lane21_data   ;

    assign reg__scntl__lane22_ready = reg__scntl__ready [22]    ;
    assign scntl__reg__valid [22]   = scntl__reg__lane22_valid  ;
    assign scntl__reg__data  [22]   = scntl__reg__lane22_data   ;

    assign reg__scntl__lane23_ready = reg__scntl__ready [23]    ;
    assign scntl__reg__valid [23]   = scntl__reg__lane23_valid  ;
    assign scntl__reg__data  [23]   = scntl__reg__lane23_data   ;

    assign reg__scntl__lane24_ready = reg__scntl__ready [24]    ;
    assign scntl__reg__valid [24]   = scntl__reg__lane24_valid  ;
    assign scntl__reg__data  [24]   = scntl__reg__lane24_data   ;

    assign reg__scntl__lane25_ready = reg__scntl__ready [25]    ;
    assign scntl__reg__valid [25]   = scntl__reg__lane25_valid  ;
    assign scntl__reg__data  [25]   = scntl__reg__lane25_data   ;

    assign reg__scntl__lane26_ready = reg__scntl__ready [26]    ;
    assign scntl__reg__valid [26]   = scntl__reg__lane26_valid  ;
    assign scntl__reg__data  [26]   = scntl__reg__lane26_data   ;

    assign reg__scntl__lane27_ready = reg__scntl__ready [27]    ;
    assign scntl__reg__valid [27]   = scntl__reg__lane27_valid  ;
    assign scntl__reg__data  [27]   = scntl__reg__lane27_data   ;

    assign reg__scntl__lane28_ready = reg__scntl__ready [28]    ;
    assign scntl__reg__valid [28]   = scntl__reg__lane28_valid  ;
    assign scntl__reg__data  [28]   = scntl__reg__lane28_data   ;

    assign reg__scntl__lane29_ready = reg__scntl__ready [29]    ;
    assign scntl__reg__valid [29]   = scntl__reg__lane29_valid  ;
    assign scntl__reg__data  [29]   = scntl__reg__lane29_data   ;

    assign reg__scntl__lane30_ready = reg__scntl__ready [30]    ;
    assign scntl__reg__valid [30]   = scntl__reg__lane30_valid  ;
    assign scntl__reg__data  [30]   = scntl__reg__lane30_data   ;

    assign reg__scntl__lane31_ready = reg__scntl__ready [31]    ;
    assign scntl__reg__valid [31]   = scntl__reg__lane31_valid  ;
    assign scntl__reg__data  [31]   = scntl__reg__lane31_data   ;

