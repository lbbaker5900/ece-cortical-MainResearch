
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe0__oob_cntl           ( DownstreamStackBusOOB[0].cb_test.std__pe__oob_cntl          ), 
        .std__pe0__oob_valid          ( DownstreamStackBusOOB[0].cb_test.std__pe__oob_valid         ), 
        .pe0__std__oob_ready          ( DownstreamStackBusOOB[0].pe__std__oob_ready                 ), 
        .std__pe0__oob_type           ( DownstreamStackBusOOB[0].cb_test.std__pe__oob_type          ), 
        .std__pe0__oob_data           ( DownstreamStackBusOOB[0].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe1__oob_cntl           ( DownstreamStackBusOOB[1].cb_test.std__pe__oob_cntl          ), 
        .std__pe1__oob_valid          ( DownstreamStackBusOOB[1].cb_test.std__pe__oob_valid         ), 
        .pe1__std__oob_ready          ( DownstreamStackBusOOB[1].pe__std__oob_ready                 ), 
        .std__pe1__oob_type           ( DownstreamStackBusOOB[1].cb_test.std__pe__oob_type          ), 
        .std__pe1__oob_data           ( DownstreamStackBusOOB[1].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe2__oob_cntl           ( DownstreamStackBusOOB[2].cb_test.std__pe__oob_cntl          ), 
        .std__pe2__oob_valid          ( DownstreamStackBusOOB[2].cb_test.std__pe__oob_valid         ), 
        .pe2__std__oob_ready          ( DownstreamStackBusOOB[2].pe__std__oob_ready                 ), 
        .std__pe2__oob_type           ( DownstreamStackBusOOB[2].cb_test.std__pe__oob_type          ), 
        .std__pe2__oob_data           ( DownstreamStackBusOOB[2].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe3__oob_cntl           ( DownstreamStackBusOOB[3].cb_test.std__pe__oob_cntl          ), 
        .std__pe3__oob_valid          ( DownstreamStackBusOOB[3].cb_test.std__pe__oob_valid         ), 
        .pe3__std__oob_ready          ( DownstreamStackBusOOB[3].pe__std__oob_ready                 ), 
        .std__pe3__oob_type           ( DownstreamStackBusOOB[3].cb_test.std__pe__oob_type          ), 
        .std__pe3__oob_data           ( DownstreamStackBusOOB[3].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe4__oob_cntl           ( DownstreamStackBusOOB[4].cb_test.std__pe__oob_cntl          ), 
        .std__pe4__oob_valid          ( DownstreamStackBusOOB[4].cb_test.std__pe__oob_valid         ), 
        .pe4__std__oob_ready          ( DownstreamStackBusOOB[4].pe__std__oob_ready                 ), 
        .std__pe4__oob_type           ( DownstreamStackBusOOB[4].cb_test.std__pe__oob_type          ), 
        .std__pe4__oob_data           ( DownstreamStackBusOOB[4].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe5__oob_cntl           ( DownstreamStackBusOOB[5].cb_test.std__pe__oob_cntl          ), 
        .std__pe5__oob_valid          ( DownstreamStackBusOOB[5].cb_test.std__pe__oob_valid         ), 
        .pe5__std__oob_ready          ( DownstreamStackBusOOB[5].pe__std__oob_ready                 ), 
        .std__pe5__oob_type           ( DownstreamStackBusOOB[5].cb_test.std__pe__oob_type          ), 
        .std__pe5__oob_data           ( DownstreamStackBusOOB[5].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe6__oob_cntl           ( DownstreamStackBusOOB[6].cb_test.std__pe__oob_cntl          ), 
        .std__pe6__oob_valid          ( DownstreamStackBusOOB[6].cb_test.std__pe__oob_valid         ), 
        .pe6__std__oob_ready          ( DownstreamStackBusOOB[6].pe__std__oob_ready                 ), 
        .std__pe6__oob_type           ( DownstreamStackBusOOB[6].cb_test.std__pe__oob_type          ), 
        .std__pe6__oob_data           ( DownstreamStackBusOOB[6].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe7__oob_cntl           ( DownstreamStackBusOOB[7].cb_test.std__pe__oob_cntl          ), 
        .std__pe7__oob_valid          ( DownstreamStackBusOOB[7].cb_test.std__pe__oob_valid         ), 
        .pe7__std__oob_ready          ( DownstreamStackBusOOB[7].pe__std__oob_ready                 ), 
        .std__pe7__oob_type           ( DownstreamStackBusOOB[7].cb_test.std__pe__oob_type          ), 
        .std__pe7__oob_data           ( DownstreamStackBusOOB[7].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe8__oob_cntl           ( DownstreamStackBusOOB[8].cb_test.std__pe__oob_cntl          ), 
        .std__pe8__oob_valid          ( DownstreamStackBusOOB[8].cb_test.std__pe__oob_valid         ), 
        .pe8__std__oob_ready          ( DownstreamStackBusOOB[8].pe__std__oob_ready                 ), 
        .std__pe8__oob_type           ( DownstreamStackBusOOB[8].cb_test.std__pe__oob_type          ), 
        .std__pe8__oob_data           ( DownstreamStackBusOOB[8].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe9__oob_cntl           ( DownstreamStackBusOOB[9].cb_test.std__pe__oob_cntl          ), 
        .std__pe9__oob_valid          ( DownstreamStackBusOOB[9].cb_test.std__pe__oob_valid         ), 
        .pe9__std__oob_ready          ( DownstreamStackBusOOB[9].pe__std__oob_ready                 ), 
        .std__pe9__oob_type           ( DownstreamStackBusOOB[9].cb_test.std__pe__oob_type          ), 
        .std__pe9__oob_data           ( DownstreamStackBusOOB[9].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe10__oob_cntl           ( DownstreamStackBusOOB[10].cb_test.std__pe__oob_cntl          ), 
        .std__pe10__oob_valid          ( DownstreamStackBusOOB[10].cb_test.std__pe__oob_valid         ), 
        .pe10__std__oob_ready          ( DownstreamStackBusOOB[10].pe__std__oob_ready                 ), 
        .std__pe10__oob_type           ( DownstreamStackBusOOB[10].cb_test.std__pe__oob_type          ), 
        .std__pe10__oob_data           ( DownstreamStackBusOOB[10].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe11__oob_cntl           ( DownstreamStackBusOOB[11].cb_test.std__pe__oob_cntl          ), 
        .std__pe11__oob_valid          ( DownstreamStackBusOOB[11].cb_test.std__pe__oob_valid         ), 
        .pe11__std__oob_ready          ( DownstreamStackBusOOB[11].pe__std__oob_ready                 ), 
        .std__pe11__oob_type           ( DownstreamStackBusOOB[11].cb_test.std__pe__oob_type          ), 
        .std__pe11__oob_data           ( DownstreamStackBusOOB[11].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe12__oob_cntl           ( DownstreamStackBusOOB[12].cb_test.std__pe__oob_cntl          ), 
        .std__pe12__oob_valid          ( DownstreamStackBusOOB[12].cb_test.std__pe__oob_valid         ), 
        .pe12__std__oob_ready          ( DownstreamStackBusOOB[12].pe__std__oob_ready                 ), 
        .std__pe12__oob_type           ( DownstreamStackBusOOB[12].cb_test.std__pe__oob_type          ), 
        .std__pe12__oob_data           ( DownstreamStackBusOOB[12].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe13__oob_cntl           ( DownstreamStackBusOOB[13].cb_test.std__pe__oob_cntl          ), 
        .std__pe13__oob_valid          ( DownstreamStackBusOOB[13].cb_test.std__pe__oob_valid         ), 
        .pe13__std__oob_ready          ( DownstreamStackBusOOB[13].pe__std__oob_ready                 ), 
        .std__pe13__oob_type           ( DownstreamStackBusOOB[13].cb_test.std__pe__oob_type          ), 
        .std__pe13__oob_data           ( DownstreamStackBusOOB[13].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe14__oob_cntl           ( DownstreamStackBusOOB[14].cb_test.std__pe__oob_cntl          ), 
        .std__pe14__oob_valid          ( DownstreamStackBusOOB[14].cb_test.std__pe__oob_valid         ), 
        .pe14__std__oob_ready          ( DownstreamStackBusOOB[14].pe__std__oob_ready                 ), 
        .std__pe14__oob_type           ( DownstreamStackBusOOB[14].cb_test.std__pe__oob_type          ), 
        .std__pe14__oob_data           ( DownstreamStackBusOOB[14].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe15__oob_cntl           ( DownstreamStackBusOOB[15].cb_test.std__pe__oob_cntl          ), 
        .std__pe15__oob_valid          ( DownstreamStackBusOOB[15].cb_test.std__pe__oob_valid         ), 
        .pe15__std__oob_ready          ( DownstreamStackBusOOB[15].pe__std__oob_ready                 ), 
        .std__pe15__oob_type           ( DownstreamStackBusOOB[15].cb_test.std__pe__oob_type          ), 
        .std__pe15__oob_data           ( DownstreamStackBusOOB[15].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe16__oob_cntl           ( DownstreamStackBusOOB[16].cb_test.std__pe__oob_cntl          ), 
        .std__pe16__oob_valid          ( DownstreamStackBusOOB[16].cb_test.std__pe__oob_valid         ), 
        .pe16__std__oob_ready          ( DownstreamStackBusOOB[16].pe__std__oob_ready                 ), 
        .std__pe16__oob_type           ( DownstreamStackBusOOB[16].cb_test.std__pe__oob_type          ), 
        .std__pe16__oob_data           ( DownstreamStackBusOOB[16].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe17__oob_cntl           ( DownstreamStackBusOOB[17].cb_test.std__pe__oob_cntl          ), 
        .std__pe17__oob_valid          ( DownstreamStackBusOOB[17].cb_test.std__pe__oob_valid         ), 
        .pe17__std__oob_ready          ( DownstreamStackBusOOB[17].pe__std__oob_ready                 ), 
        .std__pe17__oob_type           ( DownstreamStackBusOOB[17].cb_test.std__pe__oob_type          ), 
        .std__pe17__oob_data           ( DownstreamStackBusOOB[17].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe18__oob_cntl           ( DownstreamStackBusOOB[18].cb_test.std__pe__oob_cntl          ), 
        .std__pe18__oob_valid          ( DownstreamStackBusOOB[18].cb_test.std__pe__oob_valid         ), 
        .pe18__std__oob_ready          ( DownstreamStackBusOOB[18].pe__std__oob_ready                 ), 
        .std__pe18__oob_type           ( DownstreamStackBusOOB[18].cb_test.std__pe__oob_type          ), 
        .std__pe18__oob_data           ( DownstreamStackBusOOB[18].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe19__oob_cntl           ( DownstreamStackBusOOB[19].cb_test.std__pe__oob_cntl          ), 
        .std__pe19__oob_valid          ( DownstreamStackBusOOB[19].cb_test.std__pe__oob_valid         ), 
        .pe19__std__oob_ready          ( DownstreamStackBusOOB[19].pe__std__oob_ready                 ), 
        .std__pe19__oob_type           ( DownstreamStackBusOOB[19].cb_test.std__pe__oob_type          ), 
        .std__pe19__oob_data           ( DownstreamStackBusOOB[19].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe20__oob_cntl           ( DownstreamStackBusOOB[20].cb_test.std__pe__oob_cntl          ), 
        .std__pe20__oob_valid          ( DownstreamStackBusOOB[20].cb_test.std__pe__oob_valid         ), 
        .pe20__std__oob_ready          ( DownstreamStackBusOOB[20].pe__std__oob_ready                 ), 
        .std__pe20__oob_type           ( DownstreamStackBusOOB[20].cb_test.std__pe__oob_type          ), 
        .std__pe20__oob_data           ( DownstreamStackBusOOB[20].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe21__oob_cntl           ( DownstreamStackBusOOB[21].cb_test.std__pe__oob_cntl          ), 
        .std__pe21__oob_valid          ( DownstreamStackBusOOB[21].cb_test.std__pe__oob_valid         ), 
        .pe21__std__oob_ready          ( DownstreamStackBusOOB[21].pe__std__oob_ready                 ), 
        .std__pe21__oob_type           ( DownstreamStackBusOOB[21].cb_test.std__pe__oob_type          ), 
        .std__pe21__oob_data           ( DownstreamStackBusOOB[21].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe22__oob_cntl           ( DownstreamStackBusOOB[22].cb_test.std__pe__oob_cntl          ), 
        .std__pe22__oob_valid          ( DownstreamStackBusOOB[22].cb_test.std__pe__oob_valid         ), 
        .pe22__std__oob_ready          ( DownstreamStackBusOOB[22].pe__std__oob_ready                 ), 
        .std__pe22__oob_type           ( DownstreamStackBusOOB[22].cb_test.std__pe__oob_type          ), 
        .std__pe22__oob_data           ( DownstreamStackBusOOB[22].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe23__oob_cntl           ( DownstreamStackBusOOB[23].cb_test.std__pe__oob_cntl          ), 
        .std__pe23__oob_valid          ( DownstreamStackBusOOB[23].cb_test.std__pe__oob_valid         ), 
        .pe23__std__oob_ready          ( DownstreamStackBusOOB[23].pe__std__oob_ready                 ), 
        .std__pe23__oob_type           ( DownstreamStackBusOOB[23].cb_test.std__pe__oob_type          ), 
        .std__pe23__oob_data           ( DownstreamStackBusOOB[23].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe24__oob_cntl           ( DownstreamStackBusOOB[24].cb_test.std__pe__oob_cntl          ), 
        .std__pe24__oob_valid          ( DownstreamStackBusOOB[24].cb_test.std__pe__oob_valid         ), 
        .pe24__std__oob_ready          ( DownstreamStackBusOOB[24].pe__std__oob_ready                 ), 
        .std__pe24__oob_type           ( DownstreamStackBusOOB[24].cb_test.std__pe__oob_type          ), 
        .std__pe24__oob_data           ( DownstreamStackBusOOB[24].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe25__oob_cntl           ( DownstreamStackBusOOB[25].cb_test.std__pe__oob_cntl          ), 
        .std__pe25__oob_valid          ( DownstreamStackBusOOB[25].cb_test.std__pe__oob_valid         ), 
        .pe25__std__oob_ready          ( DownstreamStackBusOOB[25].pe__std__oob_ready                 ), 
        .std__pe25__oob_type           ( DownstreamStackBusOOB[25].cb_test.std__pe__oob_type          ), 
        .std__pe25__oob_data           ( DownstreamStackBusOOB[25].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe26__oob_cntl           ( DownstreamStackBusOOB[26].cb_test.std__pe__oob_cntl          ), 
        .std__pe26__oob_valid          ( DownstreamStackBusOOB[26].cb_test.std__pe__oob_valid         ), 
        .pe26__std__oob_ready          ( DownstreamStackBusOOB[26].pe__std__oob_ready                 ), 
        .std__pe26__oob_type           ( DownstreamStackBusOOB[26].cb_test.std__pe__oob_type          ), 
        .std__pe26__oob_data           ( DownstreamStackBusOOB[26].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe27__oob_cntl           ( DownstreamStackBusOOB[27].cb_test.std__pe__oob_cntl          ), 
        .std__pe27__oob_valid          ( DownstreamStackBusOOB[27].cb_test.std__pe__oob_valid         ), 
        .pe27__std__oob_ready          ( DownstreamStackBusOOB[27].pe__std__oob_ready                 ), 
        .std__pe27__oob_type           ( DownstreamStackBusOOB[27].cb_test.std__pe__oob_type          ), 
        .std__pe27__oob_data           ( DownstreamStackBusOOB[27].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe28__oob_cntl           ( DownstreamStackBusOOB[28].cb_test.std__pe__oob_cntl          ), 
        .std__pe28__oob_valid          ( DownstreamStackBusOOB[28].cb_test.std__pe__oob_valid         ), 
        .pe28__std__oob_ready          ( DownstreamStackBusOOB[28].pe__std__oob_ready                 ), 
        .std__pe28__oob_type           ( DownstreamStackBusOOB[28].cb_test.std__pe__oob_type          ), 
        .std__pe28__oob_data           ( DownstreamStackBusOOB[28].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe29__oob_cntl           ( DownstreamStackBusOOB[29].cb_test.std__pe__oob_cntl          ), 
        .std__pe29__oob_valid          ( DownstreamStackBusOOB[29].cb_test.std__pe__oob_valid         ), 
        .pe29__std__oob_ready          ( DownstreamStackBusOOB[29].pe__std__oob_ready                 ), 
        .std__pe29__oob_type           ( DownstreamStackBusOOB[29].cb_test.std__pe__oob_type          ), 
        .std__pe29__oob_data           ( DownstreamStackBusOOB[29].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe30__oob_cntl           ( DownstreamStackBusOOB[30].cb_test.std__pe__oob_cntl          ), 
        .std__pe30__oob_valid          ( DownstreamStackBusOOB[30].cb_test.std__pe__oob_valid         ), 
        .pe30__std__oob_ready          ( DownstreamStackBusOOB[30].pe__std__oob_ready                 ), 
        .std__pe30__oob_type           ( DownstreamStackBusOOB[30].cb_test.std__pe__oob_type          ), 
        .std__pe30__oob_data           ( DownstreamStackBusOOB[30].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe31__oob_cntl           ( DownstreamStackBusOOB[31].cb_test.std__pe__oob_cntl          ), 
        .std__pe31__oob_valid          ( DownstreamStackBusOOB[31].cb_test.std__pe__oob_valid         ), 
        .pe31__std__oob_ready          ( DownstreamStackBusOOB[31].pe__std__oob_ready                 ), 
        .std__pe31__oob_type           ( DownstreamStackBusOOB[31].cb_test.std__pe__oob_type          ), 
        .std__pe31__oob_data           ( DownstreamStackBusOOB[31].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe32__oob_cntl           ( DownstreamStackBusOOB[32].cb_test.std__pe__oob_cntl          ), 
        .std__pe32__oob_valid          ( DownstreamStackBusOOB[32].cb_test.std__pe__oob_valid         ), 
        .pe32__std__oob_ready          ( DownstreamStackBusOOB[32].pe__std__oob_ready                 ), 
        .std__pe32__oob_type           ( DownstreamStackBusOOB[32].cb_test.std__pe__oob_type          ), 
        .std__pe32__oob_data           ( DownstreamStackBusOOB[32].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe33__oob_cntl           ( DownstreamStackBusOOB[33].cb_test.std__pe__oob_cntl          ), 
        .std__pe33__oob_valid          ( DownstreamStackBusOOB[33].cb_test.std__pe__oob_valid         ), 
        .pe33__std__oob_ready          ( DownstreamStackBusOOB[33].pe__std__oob_ready                 ), 
        .std__pe33__oob_type           ( DownstreamStackBusOOB[33].cb_test.std__pe__oob_type          ), 
        .std__pe33__oob_data           ( DownstreamStackBusOOB[33].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe34__oob_cntl           ( DownstreamStackBusOOB[34].cb_test.std__pe__oob_cntl          ), 
        .std__pe34__oob_valid          ( DownstreamStackBusOOB[34].cb_test.std__pe__oob_valid         ), 
        .pe34__std__oob_ready          ( DownstreamStackBusOOB[34].pe__std__oob_ready                 ), 
        .std__pe34__oob_type           ( DownstreamStackBusOOB[34].cb_test.std__pe__oob_type          ), 
        .std__pe34__oob_data           ( DownstreamStackBusOOB[34].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe35__oob_cntl           ( DownstreamStackBusOOB[35].cb_test.std__pe__oob_cntl          ), 
        .std__pe35__oob_valid          ( DownstreamStackBusOOB[35].cb_test.std__pe__oob_valid         ), 
        .pe35__std__oob_ready          ( DownstreamStackBusOOB[35].pe__std__oob_ready                 ), 
        .std__pe35__oob_type           ( DownstreamStackBusOOB[35].cb_test.std__pe__oob_type          ), 
        .std__pe35__oob_data           ( DownstreamStackBusOOB[35].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe36__oob_cntl           ( DownstreamStackBusOOB[36].cb_test.std__pe__oob_cntl          ), 
        .std__pe36__oob_valid          ( DownstreamStackBusOOB[36].cb_test.std__pe__oob_valid         ), 
        .pe36__std__oob_ready          ( DownstreamStackBusOOB[36].pe__std__oob_ready                 ), 
        .std__pe36__oob_type           ( DownstreamStackBusOOB[36].cb_test.std__pe__oob_type          ), 
        .std__pe36__oob_data           ( DownstreamStackBusOOB[36].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe37__oob_cntl           ( DownstreamStackBusOOB[37].cb_test.std__pe__oob_cntl          ), 
        .std__pe37__oob_valid          ( DownstreamStackBusOOB[37].cb_test.std__pe__oob_valid         ), 
        .pe37__std__oob_ready          ( DownstreamStackBusOOB[37].pe__std__oob_ready                 ), 
        .std__pe37__oob_type           ( DownstreamStackBusOOB[37].cb_test.std__pe__oob_type          ), 
        .std__pe37__oob_data           ( DownstreamStackBusOOB[37].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe38__oob_cntl           ( DownstreamStackBusOOB[38].cb_test.std__pe__oob_cntl          ), 
        .std__pe38__oob_valid          ( DownstreamStackBusOOB[38].cb_test.std__pe__oob_valid         ), 
        .pe38__std__oob_ready          ( DownstreamStackBusOOB[38].pe__std__oob_ready                 ), 
        .std__pe38__oob_type           ( DownstreamStackBusOOB[38].cb_test.std__pe__oob_type          ), 
        .std__pe38__oob_data           ( DownstreamStackBusOOB[38].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe39__oob_cntl           ( DownstreamStackBusOOB[39].cb_test.std__pe__oob_cntl          ), 
        .std__pe39__oob_valid          ( DownstreamStackBusOOB[39].cb_test.std__pe__oob_valid         ), 
        .pe39__std__oob_ready          ( DownstreamStackBusOOB[39].pe__std__oob_ready                 ), 
        .std__pe39__oob_type           ( DownstreamStackBusOOB[39].cb_test.std__pe__oob_type          ), 
        .std__pe39__oob_data           ( DownstreamStackBusOOB[39].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe40__oob_cntl           ( DownstreamStackBusOOB[40].cb_test.std__pe__oob_cntl          ), 
        .std__pe40__oob_valid          ( DownstreamStackBusOOB[40].cb_test.std__pe__oob_valid         ), 
        .pe40__std__oob_ready          ( DownstreamStackBusOOB[40].pe__std__oob_ready                 ), 
        .std__pe40__oob_type           ( DownstreamStackBusOOB[40].cb_test.std__pe__oob_type          ), 
        .std__pe40__oob_data           ( DownstreamStackBusOOB[40].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe41__oob_cntl           ( DownstreamStackBusOOB[41].cb_test.std__pe__oob_cntl          ), 
        .std__pe41__oob_valid          ( DownstreamStackBusOOB[41].cb_test.std__pe__oob_valid         ), 
        .pe41__std__oob_ready          ( DownstreamStackBusOOB[41].pe__std__oob_ready                 ), 
        .std__pe41__oob_type           ( DownstreamStackBusOOB[41].cb_test.std__pe__oob_type          ), 
        .std__pe41__oob_data           ( DownstreamStackBusOOB[41].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe42__oob_cntl           ( DownstreamStackBusOOB[42].cb_test.std__pe__oob_cntl          ), 
        .std__pe42__oob_valid          ( DownstreamStackBusOOB[42].cb_test.std__pe__oob_valid         ), 
        .pe42__std__oob_ready          ( DownstreamStackBusOOB[42].pe__std__oob_ready                 ), 
        .std__pe42__oob_type           ( DownstreamStackBusOOB[42].cb_test.std__pe__oob_type          ), 
        .std__pe42__oob_data           ( DownstreamStackBusOOB[42].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe43__oob_cntl           ( DownstreamStackBusOOB[43].cb_test.std__pe__oob_cntl          ), 
        .std__pe43__oob_valid          ( DownstreamStackBusOOB[43].cb_test.std__pe__oob_valid         ), 
        .pe43__std__oob_ready          ( DownstreamStackBusOOB[43].pe__std__oob_ready                 ), 
        .std__pe43__oob_type           ( DownstreamStackBusOOB[43].cb_test.std__pe__oob_type          ), 
        .std__pe43__oob_data           ( DownstreamStackBusOOB[43].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe44__oob_cntl           ( DownstreamStackBusOOB[44].cb_test.std__pe__oob_cntl          ), 
        .std__pe44__oob_valid          ( DownstreamStackBusOOB[44].cb_test.std__pe__oob_valid         ), 
        .pe44__std__oob_ready          ( DownstreamStackBusOOB[44].pe__std__oob_ready                 ), 
        .std__pe44__oob_type           ( DownstreamStackBusOOB[44].cb_test.std__pe__oob_type          ), 
        .std__pe44__oob_data           ( DownstreamStackBusOOB[44].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe45__oob_cntl           ( DownstreamStackBusOOB[45].cb_test.std__pe__oob_cntl          ), 
        .std__pe45__oob_valid          ( DownstreamStackBusOOB[45].cb_test.std__pe__oob_valid         ), 
        .pe45__std__oob_ready          ( DownstreamStackBusOOB[45].pe__std__oob_ready                 ), 
        .std__pe45__oob_type           ( DownstreamStackBusOOB[45].cb_test.std__pe__oob_type          ), 
        .std__pe45__oob_data           ( DownstreamStackBusOOB[45].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe46__oob_cntl           ( DownstreamStackBusOOB[46].cb_test.std__pe__oob_cntl          ), 
        .std__pe46__oob_valid          ( DownstreamStackBusOOB[46].cb_test.std__pe__oob_valid         ), 
        .pe46__std__oob_ready          ( DownstreamStackBusOOB[46].pe__std__oob_ready                 ), 
        .std__pe46__oob_type           ( DownstreamStackBusOOB[46].cb_test.std__pe__oob_type          ), 
        .std__pe46__oob_data           ( DownstreamStackBusOOB[46].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe47__oob_cntl           ( DownstreamStackBusOOB[47].cb_test.std__pe__oob_cntl          ), 
        .std__pe47__oob_valid          ( DownstreamStackBusOOB[47].cb_test.std__pe__oob_valid         ), 
        .pe47__std__oob_ready          ( DownstreamStackBusOOB[47].pe__std__oob_ready                 ), 
        .std__pe47__oob_type           ( DownstreamStackBusOOB[47].cb_test.std__pe__oob_type          ), 
        .std__pe47__oob_data           ( DownstreamStackBusOOB[47].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe48__oob_cntl           ( DownstreamStackBusOOB[48].cb_test.std__pe__oob_cntl          ), 
        .std__pe48__oob_valid          ( DownstreamStackBusOOB[48].cb_test.std__pe__oob_valid         ), 
        .pe48__std__oob_ready          ( DownstreamStackBusOOB[48].pe__std__oob_ready                 ), 
        .std__pe48__oob_type           ( DownstreamStackBusOOB[48].cb_test.std__pe__oob_type          ), 
        .std__pe48__oob_data           ( DownstreamStackBusOOB[48].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe49__oob_cntl           ( DownstreamStackBusOOB[49].cb_test.std__pe__oob_cntl          ), 
        .std__pe49__oob_valid          ( DownstreamStackBusOOB[49].cb_test.std__pe__oob_valid         ), 
        .pe49__std__oob_ready          ( DownstreamStackBusOOB[49].pe__std__oob_ready                 ), 
        .std__pe49__oob_type           ( DownstreamStackBusOOB[49].cb_test.std__pe__oob_type          ), 
        .std__pe49__oob_data           ( DownstreamStackBusOOB[49].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe50__oob_cntl           ( DownstreamStackBusOOB[50].cb_test.std__pe__oob_cntl          ), 
        .std__pe50__oob_valid          ( DownstreamStackBusOOB[50].cb_test.std__pe__oob_valid         ), 
        .pe50__std__oob_ready          ( DownstreamStackBusOOB[50].pe__std__oob_ready                 ), 
        .std__pe50__oob_type           ( DownstreamStackBusOOB[50].cb_test.std__pe__oob_type          ), 
        .std__pe50__oob_data           ( DownstreamStackBusOOB[50].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe51__oob_cntl           ( DownstreamStackBusOOB[51].cb_test.std__pe__oob_cntl          ), 
        .std__pe51__oob_valid          ( DownstreamStackBusOOB[51].cb_test.std__pe__oob_valid         ), 
        .pe51__std__oob_ready          ( DownstreamStackBusOOB[51].pe__std__oob_ready                 ), 
        .std__pe51__oob_type           ( DownstreamStackBusOOB[51].cb_test.std__pe__oob_type          ), 
        .std__pe51__oob_data           ( DownstreamStackBusOOB[51].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe52__oob_cntl           ( DownstreamStackBusOOB[52].cb_test.std__pe__oob_cntl          ), 
        .std__pe52__oob_valid          ( DownstreamStackBusOOB[52].cb_test.std__pe__oob_valid         ), 
        .pe52__std__oob_ready          ( DownstreamStackBusOOB[52].pe__std__oob_ready                 ), 
        .std__pe52__oob_type           ( DownstreamStackBusOOB[52].cb_test.std__pe__oob_type          ), 
        .std__pe52__oob_data           ( DownstreamStackBusOOB[52].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe53__oob_cntl           ( DownstreamStackBusOOB[53].cb_test.std__pe__oob_cntl          ), 
        .std__pe53__oob_valid          ( DownstreamStackBusOOB[53].cb_test.std__pe__oob_valid         ), 
        .pe53__std__oob_ready          ( DownstreamStackBusOOB[53].pe__std__oob_ready                 ), 
        .std__pe53__oob_type           ( DownstreamStackBusOOB[53].cb_test.std__pe__oob_type          ), 
        .std__pe53__oob_data           ( DownstreamStackBusOOB[53].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe54__oob_cntl           ( DownstreamStackBusOOB[54].cb_test.std__pe__oob_cntl          ), 
        .std__pe54__oob_valid          ( DownstreamStackBusOOB[54].cb_test.std__pe__oob_valid         ), 
        .pe54__std__oob_ready          ( DownstreamStackBusOOB[54].pe__std__oob_ready                 ), 
        .std__pe54__oob_type           ( DownstreamStackBusOOB[54].cb_test.std__pe__oob_type          ), 
        .std__pe54__oob_data           ( DownstreamStackBusOOB[54].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe55__oob_cntl           ( DownstreamStackBusOOB[55].cb_test.std__pe__oob_cntl          ), 
        .std__pe55__oob_valid          ( DownstreamStackBusOOB[55].cb_test.std__pe__oob_valid         ), 
        .pe55__std__oob_ready          ( DownstreamStackBusOOB[55].pe__std__oob_ready                 ), 
        .std__pe55__oob_type           ( DownstreamStackBusOOB[55].cb_test.std__pe__oob_type          ), 
        .std__pe55__oob_data           ( DownstreamStackBusOOB[55].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe56__oob_cntl           ( DownstreamStackBusOOB[56].cb_test.std__pe__oob_cntl          ), 
        .std__pe56__oob_valid          ( DownstreamStackBusOOB[56].cb_test.std__pe__oob_valid         ), 
        .pe56__std__oob_ready          ( DownstreamStackBusOOB[56].pe__std__oob_ready                 ), 
        .std__pe56__oob_type           ( DownstreamStackBusOOB[56].cb_test.std__pe__oob_type          ), 
        .std__pe56__oob_data           ( DownstreamStackBusOOB[56].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe57__oob_cntl           ( DownstreamStackBusOOB[57].cb_test.std__pe__oob_cntl          ), 
        .std__pe57__oob_valid          ( DownstreamStackBusOOB[57].cb_test.std__pe__oob_valid         ), 
        .pe57__std__oob_ready          ( DownstreamStackBusOOB[57].pe__std__oob_ready                 ), 
        .std__pe57__oob_type           ( DownstreamStackBusOOB[57].cb_test.std__pe__oob_type          ), 
        .std__pe57__oob_data           ( DownstreamStackBusOOB[57].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe58__oob_cntl           ( DownstreamStackBusOOB[58].cb_test.std__pe__oob_cntl          ), 
        .std__pe58__oob_valid          ( DownstreamStackBusOOB[58].cb_test.std__pe__oob_valid         ), 
        .pe58__std__oob_ready          ( DownstreamStackBusOOB[58].pe__std__oob_ready                 ), 
        .std__pe58__oob_type           ( DownstreamStackBusOOB[58].cb_test.std__pe__oob_type          ), 
        .std__pe58__oob_data           ( DownstreamStackBusOOB[58].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe59__oob_cntl           ( DownstreamStackBusOOB[59].cb_test.std__pe__oob_cntl          ), 
        .std__pe59__oob_valid          ( DownstreamStackBusOOB[59].cb_test.std__pe__oob_valid         ), 
        .pe59__std__oob_ready          ( DownstreamStackBusOOB[59].pe__std__oob_ready                 ), 
        .std__pe59__oob_type           ( DownstreamStackBusOOB[59].cb_test.std__pe__oob_type          ), 
        .std__pe59__oob_data           ( DownstreamStackBusOOB[59].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe60__oob_cntl           ( DownstreamStackBusOOB[60].cb_test.std__pe__oob_cntl          ), 
        .std__pe60__oob_valid          ( DownstreamStackBusOOB[60].cb_test.std__pe__oob_valid         ), 
        .pe60__std__oob_ready          ( DownstreamStackBusOOB[60].pe__std__oob_ready                 ), 
        .std__pe60__oob_type           ( DownstreamStackBusOOB[60].cb_test.std__pe__oob_type          ), 
        .std__pe60__oob_data           ( DownstreamStackBusOOB[60].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe61__oob_cntl           ( DownstreamStackBusOOB[61].cb_test.std__pe__oob_cntl          ), 
        .std__pe61__oob_valid          ( DownstreamStackBusOOB[61].cb_test.std__pe__oob_valid         ), 
        .pe61__std__oob_ready          ( DownstreamStackBusOOB[61].pe__std__oob_ready                 ), 
        .std__pe61__oob_type           ( DownstreamStackBusOOB[61].cb_test.std__pe__oob_type          ), 
        .std__pe61__oob_data           ( DownstreamStackBusOOB[61].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe62__oob_cntl           ( DownstreamStackBusOOB[62].cb_test.std__pe__oob_cntl          ), 
        .std__pe62__oob_valid          ( DownstreamStackBusOOB[62].cb_test.std__pe__oob_valid         ), 
        .pe62__std__oob_ready          ( DownstreamStackBusOOB[62].pe__std__oob_ready                 ), 
        .std__pe62__oob_type           ( DownstreamStackBusOOB[62].cb_test.std__pe__oob_type          ), 
        .std__pe62__oob_data           ( DownstreamStackBusOOB[62].cb_test.std__pe__oob_data          ), 
  // OOB controls how the lanes are interpreted                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .std__pe63__oob_cntl           ( DownstreamStackBusOOB[63].cb_test.std__pe__oob_cntl          ), 
        .std__pe63__oob_valid          ( DownstreamStackBusOOB[63].cb_test.std__pe__oob_valid         ), 
        .pe63__std__oob_ready          ( DownstreamStackBusOOB[63].pe__std__oob_ready                 ), 
        .std__pe63__oob_type           ( DownstreamStackBusOOB[63].cb_test.std__pe__oob_type          ), 
        .std__pe63__oob_data           ( DownstreamStackBusOOB[63].cb_test.std__pe__oob_data          ), 