
`ifdef SYNTHESIS
            // Memory port 0
            memc__sram__read_address0 ,
            sram__memc__read_data0 ,
            memc__sram__write_address0 ,
            memc__sram__write_enable0 ,
            memc__sram__write_data0 ,

            // Memory port 1
            memc__sram__read_address1 ,
            sram__memc__read_data1 ,
            memc__sram__write_address1 ,
            memc__sram__write_enable1 ,
            memc__sram__write_data1 ,

            // Memory port 2
            memc__sram__read_address2 ,
            sram__memc__read_data2 ,
            memc__sram__write_address2 ,
            memc__sram__write_enable2 ,
            memc__sram__write_data2 ,

            // Memory port 3
            memc__sram__read_address3 ,
            sram__memc__read_data3 ,
            memc__sram__write_address3 ,
            memc__sram__write_enable3 ,
            memc__sram__write_data3 ,

            // Memory port 4
            memc__sram__read_address4 ,
            sram__memc__read_data4 ,
            memc__sram__write_address4 ,
            memc__sram__write_enable4 ,
            memc__sram__write_data4 ,

            // Memory port 5
            memc__sram__read_address5 ,
            sram__memc__read_data5 ,
            memc__sram__write_address5 ,
            memc__sram__write_enable5 ,
            memc__sram__write_data5 ,

            // Memory port 6
            memc__sram__read_address6 ,
            sram__memc__read_data6 ,
            memc__sram__write_address6 ,
            memc__sram__write_enable6 ,
            memc__sram__write_data6 ,

            // Memory port 7
            memc__sram__read_address7 ,
            sram__memc__read_data7 ,
            memc__sram__write_address7 ,
            memc__sram__write_enable7 ,
            memc__sram__write_data7 ,

            // Memory port 8
            memc__sram__read_address8 ,
            sram__memc__read_data8 ,
            memc__sram__write_address8 ,
            memc__sram__write_enable8 ,
            memc__sram__write_data8 ,

            // Memory port 9
            memc__sram__read_address9 ,
            sram__memc__read_data9 ,
            memc__sram__write_address9 ,
            memc__sram__write_enable9 ,
            memc__sram__write_data9 ,

            // Memory port 10
            memc__sram__read_address10 ,
            sram__memc__read_data10 ,
            memc__sram__write_address10 ,
            memc__sram__write_enable10 ,
            memc__sram__write_data10 ,

            // Memory port 11
            memc__sram__read_address11 ,
            sram__memc__read_data11 ,
            memc__sram__write_address11 ,
            memc__sram__write_enable11 ,
            memc__sram__write_data11 ,

            // Memory port 12
            memc__sram__read_address12 ,
            sram__memc__read_data12 ,
            memc__sram__write_address12 ,
            memc__sram__write_enable12 ,
            memc__sram__write_data12 ,

            // Memory port 13
            memc__sram__read_address13 ,
            sram__memc__read_data13 ,
            memc__sram__write_address13 ,
            memc__sram__write_enable13 ,
            memc__sram__write_data13 ,

            // Memory port 14
            memc__sram__read_address14 ,
            sram__memc__read_data14 ,
            memc__sram__write_address14 ,
            memc__sram__write_enable14 ,
            memc__sram__write_data14 ,

            // Memory port 15
            memc__sram__read_address15 ,
            sram__memc__read_data15 ,
            memc__sram__write_address15 ,
            memc__sram__write_enable15 ,
            memc__sram__write_data15 ,

            // Memory port 16
            memc__sram__read_address16 ,
            sram__memc__read_data16 ,
            memc__sram__write_address16 ,
            memc__sram__write_enable16 ,
            memc__sram__write_data16 ,

            // Memory port 17
            memc__sram__read_address17 ,
            sram__memc__read_data17 ,
            memc__sram__write_address17 ,
            memc__sram__write_enable17 ,
            memc__sram__write_data17 ,

            // Memory port 18
            memc__sram__read_address18 ,
            sram__memc__read_data18 ,
            memc__sram__write_address18 ,
            memc__sram__write_enable18 ,
            memc__sram__write_data18 ,

            // Memory port 19
            memc__sram__read_address19 ,
            sram__memc__read_data19 ,
            memc__sram__write_address19 ,
            memc__sram__write_enable19 ,
            memc__sram__write_data19 ,

            // Memory port 20
            memc__sram__read_address20 ,
            sram__memc__read_data20 ,
            memc__sram__write_address20 ,
            memc__sram__write_enable20 ,
            memc__sram__write_data20 ,

            // Memory port 21
            memc__sram__read_address21 ,
            sram__memc__read_data21 ,
            memc__sram__write_address21 ,
            memc__sram__write_enable21 ,
            memc__sram__write_data21 ,

            // Memory port 22
            memc__sram__read_address22 ,
            sram__memc__read_data22 ,
            memc__sram__write_address22 ,
            memc__sram__write_enable22 ,
            memc__sram__write_data22 ,

            // Memory port 23
            memc__sram__read_address23 ,
            sram__memc__read_data23 ,
            memc__sram__write_address23 ,
            memc__sram__write_enable23 ,
            memc__sram__write_data23 ,

            // Memory port 24
            memc__sram__read_address24 ,
            sram__memc__read_data24 ,
            memc__sram__write_address24 ,
            memc__sram__write_enable24 ,
            memc__sram__write_data24 ,

            // Memory port 25
            memc__sram__read_address25 ,
            sram__memc__read_data25 ,
            memc__sram__write_address25 ,
            memc__sram__write_enable25 ,
            memc__sram__write_data25 ,

            // Memory port 26
            memc__sram__read_address26 ,
            sram__memc__read_data26 ,
            memc__sram__write_address26 ,
            memc__sram__write_enable26 ,
            memc__sram__write_data26 ,

            // Memory port 27
            memc__sram__read_address27 ,
            sram__memc__read_data27 ,
            memc__sram__write_address27 ,
            memc__sram__write_enable27 ,
            memc__sram__write_data27 ,

            // Memory port 28
            memc__sram__read_address28 ,
            sram__memc__read_data28 ,
            memc__sram__write_address28 ,
            memc__sram__write_enable28 ,
            memc__sram__write_data28 ,

            // Memory port 29
            memc__sram__read_address29 ,
            sram__memc__read_data29 ,
            memc__sram__write_address29 ,
            memc__sram__write_enable29 ,
            memc__sram__write_data29 ,

            // Memory port 30
            memc__sram__read_address30 ,
            sram__memc__read_data30 ,
            memc__sram__write_address30 ,
            memc__sram__write_enable30 ,
            memc__sram__write_data30 ,

            // Memory port 31
            memc__sram__read_address31 ,
            sram__memc__read_data31 ,
            memc__sram__write_address31 ,
            memc__sram__write_enable31 ,
            memc__sram__write_data31 ,

`endif