
  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe0__oob_cntl            ;
  wire                                        std__pe0__oob_valid           ;
  wire                                        pe0__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe0__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe0__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe1__oob_cntl            ;
  wire                                        std__pe1__oob_valid           ;
  wire                                        pe1__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe1__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe1__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe2__oob_cntl            ;
  wire                                        std__pe2__oob_valid           ;
  wire                                        pe2__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe2__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe2__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe3__oob_cntl            ;
  wire                                        std__pe3__oob_valid           ;
  wire                                        pe3__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe3__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe3__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe4__oob_cntl            ;
  wire                                        std__pe4__oob_valid           ;
  wire                                        pe4__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe4__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe4__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe5__oob_cntl            ;
  wire                                        std__pe5__oob_valid           ;
  wire                                        pe5__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe5__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe5__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe6__oob_cntl            ;
  wire                                        std__pe6__oob_valid           ;
  wire                                        pe6__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe6__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe6__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe7__oob_cntl            ;
  wire                                        std__pe7__oob_valid           ;
  wire                                        pe7__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe7__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe7__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe8__oob_cntl            ;
  wire                                        std__pe8__oob_valid           ;
  wire                                        pe8__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe8__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe8__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe9__oob_cntl            ;
  wire                                        std__pe9__oob_valid           ;
  wire                                        pe9__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe9__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe9__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe10__oob_cntl            ;
  wire                                        std__pe10__oob_valid           ;
  wire                                        pe10__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe10__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe10__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe11__oob_cntl            ;
  wire                                        std__pe11__oob_valid           ;
  wire                                        pe11__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe11__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe11__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe12__oob_cntl            ;
  wire                                        std__pe12__oob_valid           ;
  wire                                        pe12__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe12__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe12__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe13__oob_cntl            ;
  wire                                        std__pe13__oob_valid           ;
  wire                                        pe13__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe13__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe13__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe14__oob_cntl            ;
  wire                                        std__pe14__oob_valid           ;
  wire                                        pe14__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe14__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe14__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe15__oob_cntl            ;
  wire                                        std__pe15__oob_valid           ;
  wire                                        pe15__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe15__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe15__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe16__oob_cntl            ;
  wire                                        std__pe16__oob_valid           ;
  wire                                        pe16__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe16__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe16__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe17__oob_cntl            ;
  wire                                        std__pe17__oob_valid           ;
  wire                                        pe17__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe17__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe17__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe18__oob_cntl            ;
  wire                                        std__pe18__oob_valid           ;
  wire                                        pe18__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe18__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe18__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe19__oob_cntl            ;
  wire                                        std__pe19__oob_valid           ;
  wire                                        pe19__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe19__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe19__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe20__oob_cntl            ;
  wire                                        std__pe20__oob_valid           ;
  wire                                        pe20__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe20__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe20__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe21__oob_cntl            ;
  wire                                        std__pe21__oob_valid           ;
  wire                                        pe21__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe21__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe21__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe22__oob_cntl            ;
  wire                                        std__pe22__oob_valid           ;
  wire                                        pe22__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe22__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe22__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe23__oob_cntl            ;
  wire                                        std__pe23__oob_valid           ;
  wire                                        pe23__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe23__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe23__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe24__oob_cntl            ;
  wire                                        std__pe24__oob_valid           ;
  wire                                        pe24__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe24__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe24__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe25__oob_cntl            ;
  wire                                        std__pe25__oob_valid           ;
  wire                                        pe25__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe25__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe25__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe26__oob_cntl            ;
  wire                                        std__pe26__oob_valid           ;
  wire                                        pe26__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe26__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe26__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe27__oob_cntl            ;
  wire                                        std__pe27__oob_valid           ;
  wire                                        pe27__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe27__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe27__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe28__oob_cntl            ;
  wire                                        std__pe28__oob_valid           ;
  wire                                        pe28__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe28__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe28__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe29__oob_cntl            ;
  wire                                        std__pe29__oob_valid           ;
  wire                                        pe29__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe29__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe29__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe30__oob_cntl            ;
  wire                                        std__pe30__oob_valid           ;
  wire                                        pe30__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe30__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe30__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe31__oob_cntl            ;
  wire                                        std__pe31__oob_valid           ;
  wire                                        pe31__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe31__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe31__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe32__oob_cntl            ;
  wire                                        std__pe32__oob_valid           ;
  wire                                        pe32__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe32__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe32__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe33__oob_cntl            ;
  wire                                        std__pe33__oob_valid           ;
  wire                                        pe33__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe33__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe33__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe34__oob_cntl            ;
  wire                                        std__pe34__oob_valid           ;
  wire                                        pe34__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe34__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe34__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe35__oob_cntl            ;
  wire                                        std__pe35__oob_valid           ;
  wire                                        pe35__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe35__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe35__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe36__oob_cntl            ;
  wire                                        std__pe36__oob_valid           ;
  wire                                        pe36__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe36__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe36__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe37__oob_cntl            ;
  wire                                        std__pe37__oob_valid           ;
  wire                                        pe37__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe37__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe37__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe38__oob_cntl            ;
  wire                                        std__pe38__oob_valid           ;
  wire                                        pe38__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe38__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe38__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe39__oob_cntl            ;
  wire                                        std__pe39__oob_valid           ;
  wire                                        pe39__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe39__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe39__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe40__oob_cntl            ;
  wire                                        std__pe40__oob_valid           ;
  wire                                        pe40__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe40__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe40__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe41__oob_cntl            ;
  wire                                        std__pe41__oob_valid           ;
  wire                                        pe41__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe41__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe41__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe42__oob_cntl            ;
  wire                                        std__pe42__oob_valid           ;
  wire                                        pe42__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe42__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe42__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe43__oob_cntl            ;
  wire                                        std__pe43__oob_valid           ;
  wire                                        pe43__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe43__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe43__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe44__oob_cntl            ;
  wire                                        std__pe44__oob_valid           ;
  wire                                        pe44__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe44__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe44__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe45__oob_cntl            ;
  wire                                        std__pe45__oob_valid           ;
  wire                                        pe45__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe45__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe45__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe46__oob_cntl            ;
  wire                                        std__pe46__oob_valid           ;
  wire                                        pe46__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe46__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe46__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe47__oob_cntl            ;
  wire                                        std__pe47__oob_valid           ;
  wire                                        pe47__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe47__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe47__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe48__oob_cntl            ;
  wire                                        std__pe48__oob_valid           ;
  wire                                        pe48__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe48__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe48__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe49__oob_cntl            ;
  wire                                        std__pe49__oob_valid           ;
  wire                                        pe49__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe49__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe49__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe50__oob_cntl            ;
  wire                                        std__pe50__oob_valid           ;
  wire                                        pe50__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe50__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe50__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe51__oob_cntl            ;
  wire                                        std__pe51__oob_valid           ;
  wire                                        pe51__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe51__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe51__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe52__oob_cntl            ;
  wire                                        std__pe52__oob_valid           ;
  wire                                        pe52__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe52__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe52__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe53__oob_cntl            ;
  wire                                        std__pe53__oob_valid           ;
  wire                                        pe53__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe53__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe53__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe54__oob_cntl            ;
  wire                                        std__pe54__oob_valid           ;
  wire                                        pe54__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe54__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe54__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe55__oob_cntl            ;
  wire                                        std__pe55__oob_valid           ;
  wire                                        pe55__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe55__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe55__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe56__oob_cntl            ;
  wire                                        std__pe56__oob_valid           ;
  wire                                        pe56__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe56__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe56__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe57__oob_cntl            ;
  wire                                        std__pe57__oob_valid           ;
  wire                                        pe57__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe57__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe57__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe58__oob_cntl            ;
  wire                                        std__pe58__oob_valid           ;
  wire                                        pe58__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe58__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe58__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe59__oob_cntl            ;
  wire                                        std__pe59__oob_valid           ;
  wire                                        pe59__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe59__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe59__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe60__oob_cntl            ;
  wire                                        std__pe60__oob_valid           ;
  wire                                        pe60__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe60__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe60__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe61__oob_cntl            ;
  wire                                        std__pe61__oob_valid           ;
  wire                                        pe61__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe61__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe61__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe62__oob_cntl            ;
  wire                                        std__pe62__oob_valid           ;
  wire                                        pe62__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe62__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe62__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe63__oob_cntl            ;
  wire                                        std__pe63__oob_valid           ;
  wire                                        pe63__std__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe63__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      std__pe63__oob_data            ;
