
  // DMA port 0 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data0       ; 
  wire                                        memc__dma__read_data_valid0 ; 

  // DMA port 1 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data1       ; 
  wire                                        memc__dma__read_data_valid1 ; 

  // DMA port 2 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data2       ; 
  wire                                        memc__dma__read_data_valid2 ; 

  // DMA port 3 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data3       ; 
  wire                                        memc__dma__read_data_valid3 ; 

  // DMA port 4 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data4       ; 
  wire                                        memc__dma__read_data_valid4 ; 

  // DMA port 5 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data5       ; 
  wire                                        memc__dma__read_data_valid5 ; 

  // DMA port 6 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data6       ; 
  wire                                        memc__dma__read_data_valid6 ; 

  // DMA port 7 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data7       ; 
  wire                                        memc__dma__read_data_valid7 ; 

  // DMA port 8 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data8       ; 
  wire                                        memc__dma__read_data_valid8 ; 

  // DMA port 9 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data9       ; 
  wire                                        memc__dma__read_data_valid9 ; 

  // DMA port 10 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data10       ; 
  wire                                        memc__dma__read_data_valid10 ; 

  // DMA port 11 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data11       ; 
  wire                                        memc__dma__read_data_valid11 ; 

  // DMA port 12 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data12       ; 
  wire                                        memc__dma__read_data_valid12 ; 

  // DMA port 13 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data13       ; 
  wire                                        memc__dma__read_data_valid13 ; 

  // DMA port 14 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data14       ; 
  wire                                        memc__dma__read_data_valid14 ; 

  // DMA port 15 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data15       ; 
  wire                                        memc__dma__read_data_valid15 ; 

  // DMA port 16 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data16       ; 
  wire                                        memc__dma__read_data_valid16 ; 

  // DMA port 17 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data17       ; 
  wire                                        memc__dma__read_data_valid17 ; 

  // DMA port 18 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data18       ; 
  wire                                        memc__dma__read_data_valid18 ; 

  // DMA port 19 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data19       ; 
  wire                                        memc__dma__read_data_valid19 ; 

  // DMA port 20 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data20       ; 
  wire                                        memc__dma__read_data_valid20 ; 

  // DMA port 21 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data21       ; 
  wire                                        memc__dma__read_data_valid21 ; 

  // DMA port 22 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data22       ; 
  wire                                        memc__dma__read_data_valid22 ; 

  // DMA port 23 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data23       ; 
  wire                                        memc__dma__read_data_valid23 ; 

  // DMA port 24 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data24       ; 
  wire                                        memc__dma__read_data_valid24 ; 

  // DMA port 25 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data25       ; 
  wire                                        memc__dma__read_data_valid25 ; 

  // DMA port 26 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data26       ; 
  wire                                        memc__dma__read_data_valid26 ; 

  // DMA port 27 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data27       ; 
  wire                                        memc__dma__read_data_valid27 ; 

  // DMA port 28 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data28       ; 
  wire                                        memc__dma__read_data_valid28 ; 

  // DMA port 29 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data29       ; 
  wire                                        memc__dma__read_data_valid29 ; 

  // DMA port 30 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data30       ; 
  wire                                        memc__dma__read_data_valid30 ; 

  // DMA port 31 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data31       ; 
  wire                                        memc__dma__read_data_valid31 ; 


  // What bank is the LDST accessing
  // Bank0
  wire ldst_write_addr_to_bank0      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire ldst_read_addr_to_bank0       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire ldst_write_request_to_bank0   =  ldst_write_addr_to_bank0    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank0    =  ldst_write_request_to_bank0 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank0    =  ldst_read_addr_to_bank0      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank0     =  ldst_read_request_to_bank0   & memc__ldst__read_ready   ;                                         
  // Bank1
  wire ldst_write_addr_to_bank1      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire ldst_read_addr_to_bank1       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire ldst_write_request_to_bank1   =  ldst_write_addr_to_bank1    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank1    =  ldst_write_request_to_bank1 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank1    =  ldst_read_addr_to_bank1      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank1     =  ldst_read_request_to_bank1   & memc__ldst__read_ready   ;                                         
  // Bank2
  wire ldst_write_addr_to_bank2      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire ldst_read_addr_to_bank2       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire ldst_write_request_to_bank2   =  ldst_write_addr_to_bank2    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank2    =  ldst_write_request_to_bank2 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank2    =  ldst_read_addr_to_bank2      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank2     =  ldst_read_request_to_bank2   & memc__ldst__read_ready   ;                                         
  // Bank3
  wire ldst_write_addr_to_bank3      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire ldst_read_addr_to_bank3       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire ldst_write_request_to_bank3   =  ldst_write_addr_to_bank3    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank3    =  ldst_write_request_to_bank3 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank3    =  ldst_read_addr_to_bank3      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank3     =  ldst_read_request_to_bank3   & memc__ldst__read_ready   ;                                         
  // Bank4
  wire ldst_write_addr_to_bank4      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire ldst_read_addr_to_bank4       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire ldst_write_request_to_bank4   =  ldst_write_addr_to_bank4    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank4    =  ldst_write_request_to_bank4 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank4    =  ldst_read_addr_to_bank4      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank4     =  ldst_read_request_to_bank4   & memc__ldst__read_ready   ;                                         
  // Bank5
  wire ldst_write_addr_to_bank5      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire ldst_read_addr_to_bank5       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire ldst_write_request_to_bank5   =  ldst_write_addr_to_bank5    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank5    =  ldst_write_request_to_bank5 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank5    =  ldst_read_addr_to_bank5      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank5     =  ldst_read_request_to_bank5   & memc__ldst__read_ready   ;                                         
  // Bank6
  wire ldst_write_addr_to_bank6      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire ldst_read_addr_to_bank6       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire ldst_write_request_to_bank6   =  ldst_write_addr_to_bank6    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank6    =  ldst_write_request_to_bank6 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank6    =  ldst_read_addr_to_bank6      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank6     =  ldst_read_request_to_bank6   & memc__ldst__read_ready   ;                                         
  // Bank7
  wire ldst_write_addr_to_bank7      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire ldst_read_addr_to_bank7       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire ldst_write_request_to_bank7   =  ldst_write_addr_to_bank7    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank7    =  ldst_write_request_to_bank7 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank7    =  ldst_read_addr_to_bank7      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank7     =  ldst_read_request_to_bank7   & memc__ldst__read_ready   ;                                         
  // Bank8
  wire ldst_write_addr_to_bank8      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire ldst_read_addr_to_bank8       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire ldst_write_request_to_bank8   =  ldst_write_addr_to_bank8    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank8    =  ldst_write_request_to_bank8 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank8    =  ldst_read_addr_to_bank8      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank8     =  ldst_read_request_to_bank8   & memc__ldst__read_ready   ;                                         
  // Bank9
  wire ldst_write_addr_to_bank9      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire ldst_read_addr_to_bank9       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire ldst_write_request_to_bank9   =  ldst_write_addr_to_bank9    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank9    =  ldst_write_request_to_bank9 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank9    =  ldst_read_addr_to_bank9      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank9     =  ldst_read_request_to_bank9   & memc__ldst__read_ready   ;                                         
  // Bank10
  wire ldst_write_addr_to_bank10      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire ldst_read_addr_to_bank10       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire ldst_write_request_to_bank10   =  ldst_write_addr_to_bank10    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank10    =  ldst_write_request_to_bank10 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank10    =  ldst_read_addr_to_bank10      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank10     =  ldst_read_request_to_bank10   & memc__ldst__read_ready   ;                                         
  // Bank11
  wire ldst_write_addr_to_bank11      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire ldst_read_addr_to_bank11       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire ldst_write_request_to_bank11   =  ldst_write_addr_to_bank11    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank11    =  ldst_write_request_to_bank11 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank11    =  ldst_read_addr_to_bank11      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank11     =  ldst_read_request_to_bank11   & memc__ldst__read_ready   ;                                         
  // Bank12
  wire ldst_write_addr_to_bank12      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire ldst_read_addr_to_bank12       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire ldst_write_request_to_bank12   =  ldst_write_addr_to_bank12    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank12    =  ldst_write_request_to_bank12 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank12    =  ldst_read_addr_to_bank12      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank12     =  ldst_read_request_to_bank12   & memc__ldst__read_ready   ;                                         
  // Bank13
  wire ldst_write_addr_to_bank13      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire ldst_read_addr_to_bank13       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire ldst_write_request_to_bank13   =  ldst_write_addr_to_bank13    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank13    =  ldst_write_request_to_bank13 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank13    =  ldst_read_addr_to_bank13      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank13     =  ldst_read_request_to_bank13   & memc__ldst__read_ready   ;                                         
  // Bank14
  wire ldst_write_addr_to_bank14      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire ldst_read_addr_to_bank14       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire ldst_write_request_to_bank14   =  ldst_write_addr_to_bank14    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank14    =  ldst_write_request_to_bank14 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank14    =  ldst_read_addr_to_bank14      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank14     =  ldst_read_request_to_bank14   & memc__ldst__read_ready   ;                                         
  // Bank15
  wire ldst_write_addr_to_bank15      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire ldst_read_addr_to_bank15       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire ldst_write_request_to_bank15   =  ldst_write_addr_to_bank15    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank15    =  ldst_write_request_to_bank15 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank15    =  ldst_read_addr_to_bank15      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank15     =  ldst_read_request_to_bank15   & memc__ldst__read_ready   ;                                         
  // Bank16
  wire ldst_write_addr_to_bank16      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire ldst_read_addr_to_bank16       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire ldst_write_request_to_bank16   =  ldst_write_addr_to_bank16    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank16    =  ldst_write_request_to_bank16 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank16    =  ldst_read_addr_to_bank16      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank16     =  ldst_read_request_to_bank16   & memc__ldst__read_ready   ;                                         
  // Bank17
  wire ldst_write_addr_to_bank17      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire ldst_read_addr_to_bank17       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire ldst_write_request_to_bank17   =  ldst_write_addr_to_bank17    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank17    =  ldst_write_request_to_bank17 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank17    =  ldst_read_addr_to_bank17      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank17     =  ldst_read_request_to_bank17   & memc__ldst__read_ready   ;                                         
  // Bank18
  wire ldst_write_addr_to_bank18      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire ldst_read_addr_to_bank18       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire ldst_write_request_to_bank18   =  ldst_write_addr_to_bank18    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank18    =  ldst_write_request_to_bank18 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank18    =  ldst_read_addr_to_bank18      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank18     =  ldst_read_request_to_bank18   & memc__ldst__read_ready   ;                                         
  // Bank19
  wire ldst_write_addr_to_bank19      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire ldst_read_addr_to_bank19       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire ldst_write_request_to_bank19   =  ldst_write_addr_to_bank19    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank19    =  ldst_write_request_to_bank19 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank19    =  ldst_read_addr_to_bank19      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank19     =  ldst_read_request_to_bank19   & memc__ldst__read_ready   ;                                         
  // Bank20
  wire ldst_write_addr_to_bank20      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire ldst_read_addr_to_bank20       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire ldst_write_request_to_bank20   =  ldst_write_addr_to_bank20    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank20    =  ldst_write_request_to_bank20 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank20    =  ldst_read_addr_to_bank20      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank20     =  ldst_read_request_to_bank20   & memc__ldst__read_ready   ;                                         
  // Bank21
  wire ldst_write_addr_to_bank21      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire ldst_read_addr_to_bank21       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire ldst_write_request_to_bank21   =  ldst_write_addr_to_bank21    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank21    =  ldst_write_request_to_bank21 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank21    =  ldst_read_addr_to_bank21      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank21     =  ldst_read_request_to_bank21   & memc__ldst__read_ready   ;                                         
  // Bank22
  wire ldst_write_addr_to_bank22      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire ldst_read_addr_to_bank22       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire ldst_write_request_to_bank22   =  ldst_write_addr_to_bank22    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank22    =  ldst_write_request_to_bank22 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank22    =  ldst_read_addr_to_bank22      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank22     =  ldst_read_request_to_bank22   & memc__ldst__read_ready   ;                                         
  // Bank23
  wire ldst_write_addr_to_bank23      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire ldst_read_addr_to_bank23       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire ldst_write_request_to_bank23   =  ldst_write_addr_to_bank23    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank23    =  ldst_write_request_to_bank23 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank23    =  ldst_read_addr_to_bank23      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank23     =  ldst_read_request_to_bank23   & memc__ldst__read_ready   ;                                         
  // Bank24
  wire ldst_write_addr_to_bank24      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire ldst_read_addr_to_bank24       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire ldst_write_request_to_bank24   =  ldst_write_addr_to_bank24    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank24    =  ldst_write_request_to_bank24 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank24    =  ldst_read_addr_to_bank24      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank24     =  ldst_read_request_to_bank24   & memc__ldst__read_ready   ;                                         
  // Bank25
  wire ldst_write_addr_to_bank25      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire ldst_read_addr_to_bank25       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire ldst_write_request_to_bank25   =  ldst_write_addr_to_bank25    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank25    =  ldst_write_request_to_bank25 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank25    =  ldst_read_addr_to_bank25      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank25     =  ldst_read_request_to_bank25   & memc__ldst__read_ready   ;                                         
  // Bank26
  wire ldst_write_addr_to_bank26      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire ldst_read_addr_to_bank26       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire ldst_write_request_to_bank26   =  ldst_write_addr_to_bank26    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank26    =  ldst_write_request_to_bank26 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank26    =  ldst_read_addr_to_bank26      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank26     =  ldst_read_request_to_bank26   & memc__ldst__read_ready   ;                                         
  // Bank27
  wire ldst_write_addr_to_bank27      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire ldst_read_addr_to_bank27       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire ldst_write_request_to_bank27   =  ldst_write_addr_to_bank27    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank27    =  ldst_write_request_to_bank27 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank27    =  ldst_read_addr_to_bank27      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank27     =  ldst_read_request_to_bank27   & memc__ldst__read_ready   ;                                         
  // Bank28
  wire ldst_write_addr_to_bank28      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire ldst_read_addr_to_bank28       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire ldst_write_request_to_bank28   =  ldst_write_addr_to_bank28    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank28    =  ldst_write_request_to_bank28 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank28    =  ldst_read_addr_to_bank28      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank28     =  ldst_read_request_to_bank28   & memc__ldst__read_ready   ;                                         
  // Bank29
  wire ldst_write_addr_to_bank29      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire ldst_read_addr_to_bank29       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire ldst_write_request_to_bank29   =  ldst_write_addr_to_bank29    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank29    =  ldst_write_request_to_bank29 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank29    =  ldst_read_addr_to_bank29      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank29     =  ldst_read_request_to_bank29   & memc__ldst__read_ready   ;                                         
  // Bank30
  wire ldst_write_addr_to_bank30      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire ldst_read_addr_to_bank30       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire ldst_write_request_to_bank30   =  ldst_write_addr_to_bank30    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank30    =  ldst_write_request_to_bank30 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank30    =  ldst_read_addr_to_bank30      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank30     =  ldst_read_request_to_bank30   & memc__ldst__read_ready   ;                                         
  // Bank31
  wire ldst_write_addr_to_bank31      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire ldst_read_addr_to_bank31       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire ldst_write_request_to_bank31   =  ldst_write_addr_to_bank31    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank31    =  ldst_write_request_to_bank31 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank31    =  ldst_read_addr_to_bank31      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank31     =  ldst_read_request_to_bank31   & memc__ldst__read_ready   ;                                         

  // What banks are the DMA's accessing
  // DMA 0
  wire read_pause0     =  dma__memc__read_pause0   ;  
  // DMA 0, bank0
  wire dma_write_addr0_to_bank0      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr0_to_bank0       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank0   =  dma_write_addr0_to_bank0  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank0    =  write_request0_to_bank0   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank0    =  dma_read_addr0_to_bank0   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank0     =  read_request0_to_bank0    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank1
  wire dma_write_addr0_to_bank1      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr0_to_bank1       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank1   =  dma_write_addr0_to_bank1  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank1    =  write_request0_to_bank1   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank1    =  dma_read_addr0_to_bank1   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank1     =  read_request0_to_bank1    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank2
  wire dma_write_addr0_to_bank2      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr0_to_bank2       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank2   =  dma_write_addr0_to_bank2  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank2    =  write_request0_to_bank2   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank2    =  dma_read_addr0_to_bank2   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank2     =  read_request0_to_bank2    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank3
  wire dma_write_addr0_to_bank3      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr0_to_bank3       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank3   =  dma_write_addr0_to_bank3  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank3    =  write_request0_to_bank3   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank3    =  dma_read_addr0_to_bank3   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank3     =  read_request0_to_bank3    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank4
  wire dma_write_addr0_to_bank4      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr0_to_bank4       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank4   =  dma_write_addr0_to_bank4  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank4    =  write_request0_to_bank4   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank4    =  dma_read_addr0_to_bank4   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank4     =  read_request0_to_bank4    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank5
  wire dma_write_addr0_to_bank5      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr0_to_bank5       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank5   =  dma_write_addr0_to_bank5  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank5    =  write_request0_to_bank5   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank5    =  dma_read_addr0_to_bank5   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank5     =  read_request0_to_bank5    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank6
  wire dma_write_addr0_to_bank6      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr0_to_bank6       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank6   =  dma_write_addr0_to_bank6  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank6    =  write_request0_to_bank6   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank6    =  dma_read_addr0_to_bank6   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank6     =  read_request0_to_bank6    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank7
  wire dma_write_addr0_to_bank7      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr0_to_bank7       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank7   =  dma_write_addr0_to_bank7  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank7    =  write_request0_to_bank7   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank7    =  dma_read_addr0_to_bank7   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank7     =  read_request0_to_bank7    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank8
  wire dma_write_addr0_to_bank8      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr0_to_bank8       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank8   =  dma_write_addr0_to_bank8  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank8    =  write_request0_to_bank8   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank8    =  dma_read_addr0_to_bank8   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank8     =  read_request0_to_bank8    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank9
  wire dma_write_addr0_to_bank9      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr0_to_bank9       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank9   =  dma_write_addr0_to_bank9  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank9    =  write_request0_to_bank9   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank9    =  dma_read_addr0_to_bank9   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank9     =  read_request0_to_bank9    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank10
  wire dma_write_addr0_to_bank10      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr0_to_bank10       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank10   =  dma_write_addr0_to_bank10  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank10    =  write_request0_to_bank10   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank10    =  dma_read_addr0_to_bank10   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank10     =  read_request0_to_bank10    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank11
  wire dma_write_addr0_to_bank11      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr0_to_bank11       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank11   =  dma_write_addr0_to_bank11  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank11    =  write_request0_to_bank11   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank11    =  dma_read_addr0_to_bank11   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank11     =  read_request0_to_bank11    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank12
  wire dma_write_addr0_to_bank12      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr0_to_bank12       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank12   =  dma_write_addr0_to_bank12  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank12    =  write_request0_to_bank12   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank12    =  dma_read_addr0_to_bank12   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank12     =  read_request0_to_bank12    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank13
  wire dma_write_addr0_to_bank13      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr0_to_bank13       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank13   =  dma_write_addr0_to_bank13  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank13    =  write_request0_to_bank13   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank13    =  dma_read_addr0_to_bank13   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank13     =  read_request0_to_bank13    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank14
  wire dma_write_addr0_to_bank14      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr0_to_bank14       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank14   =  dma_write_addr0_to_bank14  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank14    =  write_request0_to_bank14   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank14    =  dma_read_addr0_to_bank14   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank14     =  read_request0_to_bank14    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank15
  wire dma_write_addr0_to_bank15      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr0_to_bank15       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank15   =  dma_write_addr0_to_bank15  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank15    =  write_request0_to_bank15   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank15    =  dma_read_addr0_to_bank15   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank15     =  read_request0_to_bank15    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank16
  wire dma_write_addr0_to_bank16      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr0_to_bank16       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank16   =  dma_write_addr0_to_bank16  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank16    =  write_request0_to_bank16   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank16    =  dma_read_addr0_to_bank16   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank16     =  read_request0_to_bank16    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank17
  wire dma_write_addr0_to_bank17      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr0_to_bank17       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank17   =  dma_write_addr0_to_bank17  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank17    =  write_request0_to_bank17   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank17    =  dma_read_addr0_to_bank17   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank17     =  read_request0_to_bank17    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank18
  wire dma_write_addr0_to_bank18      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr0_to_bank18       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank18   =  dma_write_addr0_to_bank18  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank18    =  write_request0_to_bank18   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank18    =  dma_read_addr0_to_bank18   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank18     =  read_request0_to_bank18    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank19
  wire dma_write_addr0_to_bank19      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr0_to_bank19       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank19   =  dma_write_addr0_to_bank19  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank19    =  write_request0_to_bank19   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank19    =  dma_read_addr0_to_bank19   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank19     =  read_request0_to_bank19    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank20
  wire dma_write_addr0_to_bank20      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr0_to_bank20       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank20   =  dma_write_addr0_to_bank20  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank20    =  write_request0_to_bank20   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank20    =  dma_read_addr0_to_bank20   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank20     =  read_request0_to_bank20    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank21
  wire dma_write_addr0_to_bank21      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr0_to_bank21       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank21   =  dma_write_addr0_to_bank21  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank21    =  write_request0_to_bank21   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank21    =  dma_read_addr0_to_bank21   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank21     =  read_request0_to_bank21    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank22
  wire dma_write_addr0_to_bank22      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr0_to_bank22       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank22   =  dma_write_addr0_to_bank22  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank22    =  write_request0_to_bank22   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank22    =  dma_read_addr0_to_bank22   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank22     =  read_request0_to_bank22    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank23
  wire dma_write_addr0_to_bank23      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr0_to_bank23       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank23   =  dma_write_addr0_to_bank23  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank23    =  write_request0_to_bank23   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank23    =  dma_read_addr0_to_bank23   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank23     =  read_request0_to_bank23    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank24
  wire dma_write_addr0_to_bank24      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr0_to_bank24       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank24   =  dma_write_addr0_to_bank24  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank24    =  write_request0_to_bank24   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank24    =  dma_read_addr0_to_bank24   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank24     =  read_request0_to_bank24    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank25
  wire dma_write_addr0_to_bank25      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr0_to_bank25       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank25   =  dma_write_addr0_to_bank25  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank25    =  write_request0_to_bank25   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank25    =  dma_read_addr0_to_bank25   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank25     =  read_request0_to_bank25    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank26
  wire dma_write_addr0_to_bank26      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr0_to_bank26       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank26   =  dma_write_addr0_to_bank26  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank26    =  write_request0_to_bank26   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank26    =  dma_read_addr0_to_bank26   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank26     =  read_request0_to_bank26    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank27
  wire dma_write_addr0_to_bank27      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr0_to_bank27       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank27   =  dma_write_addr0_to_bank27  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank27    =  write_request0_to_bank27   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank27    =  dma_read_addr0_to_bank27   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank27     =  read_request0_to_bank27    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank28
  wire dma_write_addr0_to_bank28      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr0_to_bank28       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank28   =  dma_write_addr0_to_bank28  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank28    =  write_request0_to_bank28   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank28    =  dma_read_addr0_to_bank28   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank28     =  read_request0_to_bank28    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank29
  wire dma_write_addr0_to_bank29      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr0_to_bank29       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank29   =  dma_write_addr0_to_bank29  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank29    =  write_request0_to_bank29   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank29    =  dma_read_addr0_to_bank29   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank29     =  read_request0_to_bank29    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank30
  wire dma_write_addr0_to_bank30      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr0_to_bank30       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank30   =  dma_write_addr0_to_bank30  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank30    =  write_request0_to_bank30   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank30    =  dma_read_addr0_to_bank30   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank30     =  read_request0_to_bank30    & memc__dma__read_ready0   ;                                         
  // DMA 0, bank31
  wire dma_write_addr0_to_bank31      =  (dma__memc__write_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr0_to_bank31       =  (dma__memc__read_address0[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank31   =  dma_write_addr0_to_bank31  & dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank31    =  write_request0_to_bank31   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank31    =  dma_read_addr0_to_bank31   & dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank31     =  read_request0_to_bank31    & memc__dma__read_ready0   ;                                         
  // DMA 1
  wire read_pause1     =  dma__memc__read_pause1   ;  
  // DMA 1, bank0
  wire dma_write_addr1_to_bank0      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr1_to_bank0       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank0   =  dma_write_addr1_to_bank0  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank0    =  write_request1_to_bank0   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank0    =  dma_read_addr1_to_bank0   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank0     =  read_request1_to_bank0    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank1
  wire dma_write_addr1_to_bank1      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr1_to_bank1       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank1   =  dma_write_addr1_to_bank1  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank1    =  write_request1_to_bank1   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank1    =  dma_read_addr1_to_bank1   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank1     =  read_request1_to_bank1    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank2
  wire dma_write_addr1_to_bank2      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr1_to_bank2       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank2   =  dma_write_addr1_to_bank2  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank2    =  write_request1_to_bank2   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank2    =  dma_read_addr1_to_bank2   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank2     =  read_request1_to_bank2    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank3
  wire dma_write_addr1_to_bank3      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr1_to_bank3       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank3   =  dma_write_addr1_to_bank3  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank3    =  write_request1_to_bank3   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank3    =  dma_read_addr1_to_bank3   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank3     =  read_request1_to_bank3    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank4
  wire dma_write_addr1_to_bank4      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr1_to_bank4       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank4   =  dma_write_addr1_to_bank4  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank4    =  write_request1_to_bank4   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank4    =  dma_read_addr1_to_bank4   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank4     =  read_request1_to_bank4    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank5
  wire dma_write_addr1_to_bank5      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr1_to_bank5       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank5   =  dma_write_addr1_to_bank5  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank5    =  write_request1_to_bank5   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank5    =  dma_read_addr1_to_bank5   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank5     =  read_request1_to_bank5    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank6
  wire dma_write_addr1_to_bank6      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr1_to_bank6       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank6   =  dma_write_addr1_to_bank6  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank6    =  write_request1_to_bank6   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank6    =  dma_read_addr1_to_bank6   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank6     =  read_request1_to_bank6    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank7
  wire dma_write_addr1_to_bank7      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr1_to_bank7       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank7   =  dma_write_addr1_to_bank7  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank7    =  write_request1_to_bank7   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank7    =  dma_read_addr1_to_bank7   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank7     =  read_request1_to_bank7    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank8
  wire dma_write_addr1_to_bank8      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr1_to_bank8       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank8   =  dma_write_addr1_to_bank8  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank8    =  write_request1_to_bank8   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank8    =  dma_read_addr1_to_bank8   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank8     =  read_request1_to_bank8    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank9
  wire dma_write_addr1_to_bank9      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr1_to_bank9       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank9   =  dma_write_addr1_to_bank9  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank9    =  write_request1_to_bank9   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank9    =  dma_read_addr1_to_bank9   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank9     =  read_request1_to_bank9    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank10
  wire dma_write_addr1_to_bank10      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr1_to_bank10       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank10   =  dma_write_addr1_to_bank10  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank10    =  write_request1_to_bank10   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank10    =  dma_read_addr1_to_bank10   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank10     =  read_request1_to_bank10    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank11
  wire dma_write_addr1_to_bank11      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr1_to_bank11       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank11   =  dma_write_addr1_to_bank11  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank11    =  write_request1_to_bank11   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank11    =  dma_read_addr1_to_bank11   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank11     =  read_request1_to_bank11    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank12
  wire dma_write_addr1_to_bank12      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr1_to_bank12       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank12   =  dma_write_addr1_to_bank12  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank12    =  write_request1_to_bank12   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank12    =  dma_read_addr1_to_bank12   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank12     =  read_request1_to_bank12    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank13
  wire dma_write_addr1_to_bank13      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr1_to_bank13       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank13   =  dma_write_addr1_to_bank13  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank13    =  write_request1_to_bank13   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank13    =  dma_read_addr1_to_bank13   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank13     =  read_request1_to_bank13    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank14
  wire dma_write_addr1_to_bank14      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr1_to_bank14       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank14   =  dma_write_addr1_to_bank14  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank14    =  write_request1_to_bank14   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank14    =  dma_read_addr1_to_bank14   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank14     =  read_request1_to_bank14    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank15
  wire dma_write_addr1_to_bank15      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr1_to_bank15       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank15   =  dma_write_addr1_to_bank15  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank15    =  write_request1_to_bank15   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank15    =  dma_read_addr1_to_bank15   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank15     =  read_request1_to_bank15    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank16
  wire dma_write_addr1_to_bank16      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr1_to_bank16       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank16   =  dma_write_addr1_to_bank16  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank16    =  write_request1_to_bank16   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank16    =  dma_read_addr1_to_bank16   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank16     =  read_request1_to_bank16    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank17
  wire dma_write_addr1_to_bank17      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr1_to_bank17       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank17   =  dma_write_addr1_to_bank17  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank17    =  write_request1_to_bank17   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank17    =  dma_read_addr1_to_bank17   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank17     =  read_request1_to_bank17    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank18
  wire dma_write_addr1_to_bank18      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr1_to_bank18       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank18   =  dma_write_addr1_to_bank18  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank18    =  write_request1_to_bank18   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank18    =  dma_read_addr1_to_bank18   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank18     =  read_request1_to_bank18    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank19
  wire dma_write_addr1_to_bank19      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr1_to_bank19       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank19   =  dma_write_addr1_to_bank19  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank19    =  write_request1_to_bank19   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank19    =  dma_read_addr1_to_bank19   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank19     =  read_request1_to_bank19    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank20
  wire dma_write_addr1_to_bank20      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr1_to_bank20       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank20   =  dma_write_addr1_to_bank20  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank20    =  write_request1_to_bank20   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank20    =  dma_read_addr1_to_bank20   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank20     =  read_request1_to_bank20    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank21
  wire dma_write_addr1_to_bank21      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr1_to_bank21       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank21   =  dma_write_addr1_to_bank21  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank21    =  write_request1_to_bank21   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank21    =  dma_read_addr1_to_bank21   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank21     =  read_request1_to_bank21    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank22
  wire dma_write_addr1_to_bank22      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr1_to_bank22       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank22   =  dma_write_addr1_to_bank22  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank22    =  write_request1_to_bank22   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank22    =  dma_read_addr1_to_bank22   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank22     =  read_request1_to_bank22    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank23
  wire dma_write_addr1_to_bank23      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr1_to_bank23       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank23   =  dma_write_addr1_to_bank23  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank23    =  write_request1_to_bank23   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank23    =  dma_read_addr1_to_bank23   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank23     =  read_request1_to_bank23    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank24
  wire dma_write_addr1_to_bank24      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr1_to_bank24       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank24   =  dma_write_addr1_to_bank24  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank24    =  write_request1_to_bank24   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank24    =  dma_read_addr1_to_bank24   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank24     =  read_request1_to_bank24    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank25
  wire dma_write_addr1_to_bank25      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr1_to_bank25       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank25   =  dma_write_addr1_to_bank25  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank25    =  write_request1_to_bank25   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank25    =  dma_read_addr1_to_bank25   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank25     =  read_request1_to_bank25    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank26
  wire dma_write_addr1_to_bank26      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr1_to_bank26       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank26   =  dma_write_addr1_to_bank26  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank26    =  write_request1_to_bank26   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank26    =  dma_read_addr1_to_bank26   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank26     =  read_request1_to_bank26    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank27
  wire dma_write_addr1_to_bank27      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr1_to_bank27       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank27   =  dma_write_addr1_to_bank27  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank27    =  write_request1_to_bank27   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank27    =  dma_read_addr1_to_bank27   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank27     =  read_request1_to_bank27    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank28
  wire dma_write_addr1_to_bank28      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr1_to_bank28       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank28   =  dma_write_addr1_to_bank28  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank28    =  write_request1_to_bank28   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank28    =  dma_read_addr1_to_bank28   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank28     =  read_request1_to_bank28    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank29
  wire dma_write_addr1_to_bank29      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr1_to_bank29       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank29   =  dma_write_addr1_to_bank29  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank29    =  write_request1_to_bank29   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank29    =  dma_read_addr1_to_bank29   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank29     =  read_request1_to_bank29    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank30
  wire dma_write_addr1_to_bank30      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr1_to_bank30       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank30   =  dma_write_addr1_to_bank30  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank30    =  write_request1_to_bank30   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank30    =  dma_read_addr1_to_bank30   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank30     =  read_request1_to_bank30    & memc__dma__read_ready1   ;                                         
  // DMA 1, bank31
  wire dma_write_addr1_to_bank31      =  (dma__memc__write_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr1_to_bank31       =  (dma__memc__read_address1[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank31   =  dma_write_addr1_to_bank31  & dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank31    =  write_request1_to_bank31   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank31    =  dma_read_addr1_to_bank31   & dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank31     =  read_request1_to_bank31    & memc__dma__read_ready1   ;                                         
  // DMA 2
  wire read_pause2     =  dma__memc__read_pause2   ;  
  // DMA 2, bank0
  wire dma_write_addr2_to_bank0      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr2_to_bank0       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank0   =  dma_write_addr2_to_bank0  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank0    =  write_request2_to_bank0   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank0    =  dma_read_addr2_to_bank0   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank0     =  read_request2_to_bank0    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank1
  wire dma_write_addr2_to_bank1      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr2_to_bank1       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank1   =  dma_write_addr2_to_bank1  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank1    =  write_request2_to_bank1   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank1    =  dma_read_addr2_to_bank1   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank1     =  read_request2_to_bank1    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank2
  wire dma_write_addr2_to_bank2      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr2_to_bank2       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank2   =  dma_write_addr2_to_bank2  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank2    =  write_request2_to_bank2   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank2    =  dma_read_addr2_to_bank2   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank2     =  read_request2_to_bank2    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank3
  wire dma_write_addr2_to_bank3      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr2_to_bank3       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank3   =  dma_write_addr2_to_bank3  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank3    =  write_request2_to_bank3   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank3    =  dma_read_addr2_to_bank3   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank3     =  read_request2_to_bank3    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank4
  wire dma_write_addr2_to_bank4      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr2_to_bank4       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank4   =  dma_write_addr2_to_bank4  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank4    =  write_request2_to_bank4   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank4    =  dma_read_addr2_to_bank4   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank4     =  read_request2_to_bank4    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank5
  wire dma_write_addr2_to_bank5      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr2_to_bank5       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank5   =  dma_write_addr2_to_bank5  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank5    =  write_request2_to_bank5   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank5    =  dma_read_addr2_to_bank5   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank5     =  read_request2_to_bank5    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank6
  wire dma_write_addr2_to_bank6      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr2_to_bank6       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank6   =  dma_write_addr2_to_bank6  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank6    =  write_request2_to_bank6   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank6    =  dma_read_addr2_to_bank6   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank6     =  read_request2_to_bank6    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank7
  wire dma_write_addr2_to_bank7      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr2_to_bank7       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank7   =  dma_write_addr2_to_bank7  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank7    =  write_request2_to_bank7   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank7    =  dma_read_addr2_to_bank7   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank7     =  read_request2_to_bank7    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank8
  wire dma_write_addr2_to_bank8      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr2_to_bank8       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank8   =  dma_write_addr2_to_bank8  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank8    =  write_request2_to_bank8   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank8    =  dma_read_addr2_to_bank8   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank8     =  read_request2_to_bank8    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank9
  wire dma_write_addr2_to_bank9      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr2_to_bank9       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank9   =  dma_write_addr2_to_bank9  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank9    =  write_request2_to_bank9   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank9    =  dma_read_addr2_to_bank9   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank9     =  read_request2_to_bank9    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank10
  wire dma_write_addr2_to_bank10      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr2_to_bank10       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank10   =  dma_write_addr2_to_bank10  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank10    =  write_request2_to_bank10   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank10    =  dma_read_addr2_to_bank10   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank10     =  read_request2_to_bank10    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank11
  wire dma_write_addr2_to_bank11      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr2_to_bank11       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank11   =  dma_write_addr2_to_bank11  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank11    =  write_request2_to_bank11   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank11    =  dma_read_addr2_to_bank11   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank11     =  read_request2_to_bank11    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank12
  wire dma_write_addr2_to_bank12      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr2_to_bank12       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank12   =  dma_write_addr2_to_bank12  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank12    =  write_request2_to_bank12   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank12    =  dma_read_addr2_to_bank12   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank12     =  read_request2_to_bank12    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank13
  wire dma_write_addr2_to_bank13      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr2_to_bank13       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank13   =  dma_write_addr2_to_bank13  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank13    =  write_request2_to_bank13   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank13    =  dma_read_addr2_to_bank13   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank13     =  read_request2_to_bank13    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank14
  wire dma_write_addr2_to_bank14      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr2_to_bank14       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank14   =  dma_write_addr2_to_bank14  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank14    =  write_request2_to_bank14   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank14    =  dma_read_addr2_to_bank14   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank14     =  read_request2_to_bank14    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank15
  wire dma_write_addr2_to_bank15      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr2_to_bank15       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank15   =  dma_write_addr2_to_bank15  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank15    =  write_request2_to_bank15   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank15    =  dma_read_addr2_to_bank15   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank15     =  read_request2_to_bank15    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank16
  wire dma_write_addr2_to_bank16      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr2_to_bank16       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank16   =  dma_write_addr2_to_bank16  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank16    =  write_request2_to_bank16   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank16    =  dma_read_addr2_to_bank16   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank16     =  read_request2_to_bank16    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank17
  wire dma_write_addr2_to_bank17      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr2_to_bank17       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank17   =  dma_write_addr2_to_bank17  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank17    =  write_request2_to_bank17   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank17    =  dma_read_addr2_to_bank17   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank17     =  read_request2_to_bank17    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank18
  wire dma_write_addr2_to_bank18      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr2_to_bank18       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank18   =  dma_write_addr2_to_bank18  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank18    =  write_request2_to_bank18   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank18    =  dma_read_addr2_to_bank18   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank18     =  read_request2_to_bank18    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank19
  wire dma_write_addr2_to_bank19      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr2_to_bank19       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank19   =  dma_write_addr2_to_bank19  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank19    =  write_request2_to_bank19   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank19    =  dma_read_addr2_to_bank19   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank19     =  read_request2_to_bank19    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank20
  wire dma_write_addr2_to_bank20      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr2_to_bank20       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank20   =  dma_write_addr2_to_bank20  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank20    =  write_request2_to_bank20   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank20    =  dma_read_addr2_to_bank20   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank20     =  read_request2_to_bank20    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank21
  wire dma_write_addr2_to_bank21      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr2_to_bank21       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank21   =  dma_write_addr2_to_bank21  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank21    =  write_request2_to_bank21   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank21    =  dma_read_addr2_to_bank21   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank21     =  read_request2_to_bank21    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank22
  wire dma_write_addr2_to_bank22      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr2_to_bank22       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank22   =  dma_write_addr2_to_bank22  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank22    =  write_request2_to_bank22   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank22    =  dma_read_addr2_to_bank22   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank22     =  read_request2_to_bank22    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank23
  wire dma_write_addr2_to_bank23      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr2_to_bank23       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank23   =  dma_write_addr2_to_bank23  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank23    =  write_request2_to_bank23   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank23    =  dma_read_addr2_to_bank23   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank23     =  read_request2_to_bank23    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank24
  wire dma_write_addr2_to_bank24      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr2_to_bank24       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank24   =  dma_write_addr2_to_bank24  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank24    =  write_request2_to_bank24   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank24    =  dma_read_addr2_to_bank24   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank24     =  read_request2_to_bank24    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank25
  wire dma_write_addr2_to_bank25      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr2_to_bank25       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank25   =  dma_write_addr2_to_bank25  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank25    =  write_request2_to_bank25   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank25    =  dma_read_addr2_to_bank25   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank25     =  read_request2_to_bank25    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank26
  wire dma_write_addr2_to_bank26      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr2_to_bank26       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank26   =  dma_write_addr2_to_bank26  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank26    =  write_request2_to_bank26   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank26    =  dma_read_addr2_to_bank26   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank26     =  read_request2_to_bank26    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank27
  wire dma_write_addr2_to_bank27      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr2_to_bank27       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank27   =  dma_write_addr2_to_bank27  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank27    =  write_request2_to_bank27   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank27    =  dma_read_addr2_to_bank27   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank27     =  read_request2_to_bank27    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank28
  wire dma_write_addr2_to_bank28      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr2_to_bank28       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank28   =  dma_write_addr2_to_bank28  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank28    =  write_request2_to_bank28   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank28    =  dma_read_addr2_to_bank28   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank28     =  read_request2_to_bank28    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank29
  wire dma_write_addr2_to_bank29      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr2_to_bank29       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank29   =  dma_write_addr2_to_bank29  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank29    =  write_request2_to_bank29   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank29    =  dma_read_addr2_to_bank29   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank29     =  read_request2_to_bank29    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank30
  wire dma_write_addr2_to_bank30      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr2_to_bank30       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank30   =  dma_write_addr2_to_bank30  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank30    =  write_request2_to_bank30   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank30    =  dma_read_addr2_to_bank30   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank30     =  read_request2_to_bank30    & memc__dma__read_ready2   ;                                         
  // DMA 2, bank31
  wire dma_write_addr2_to_bank31      =  (dma__memc__write_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr2_to_bank31       =  (dma__memc__read_address2[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank31   =  dma_write_addr2_to_bank31  & dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank31    =  write_request2_to_bank31   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank31    =  dma_read_addr2_to_bank31   & dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank31     =  read_request2_to_bank31    & memc__dma__read_ready2   ;                                         
  // DMA 3
  wire read_pause3     =  dma__memc__read_pause3   ;  
  // DMA 3, bank0
  wire dma_write_addr3_to_bank0      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr3_to_bank0       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank0   =  dma_write_addr3_to_bank0  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank0    =  write_request3_to_bank0   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank0    =  dma_read_addr3_to_bank0   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank0     =  read_request3_to_bank0    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank1
  wire dma_write_addr3_to_bank1      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr3_to_bank1       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank1   =  dma_write_addr3_to_bank1  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank1    =  write_request3_to_bank1   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank1    =  dma_read_addr3_to_bank1   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank1     =  read_request3_to_bank1    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank2
  wire dma_write_addr3_to_bank2      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr3_to_bank2       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank2   =  dma_write_addr3_to_bank2  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank2    =  write_request3_to_bank2   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank2    =  dma_read_addr3_to_bank2   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank2     =  read_request3_to_bank2    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank3
  wire dma_write_addr3_to_bank3      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr3_to_bank3       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank3   =  dma_write_addr3_to_bank3  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank3    =  write_request3_to_bank3   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank3    =  dma_read_addr3_to_bank3   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank3     =  read_request3_to_bank3    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank4
  wire dma_write_addr3_to_bank4      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr3_to_bank4       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank4   =  dma_write_addr3_to_bank4  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank4    =  write_request3_to_bank4   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank4    =  dma_read_addr3_to_bank4   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank4     =  read_request3_to_bank4    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank5
  wire dma_write_addr3_to_bank5      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr3_to_bank5       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank5   =  dma_write_addr3_to_bank5  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank5    =  write_request3_to_bank5   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank5    =  dma_read_addr3_to_bank5   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank5     =  read_request3_to_bank5    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank6
  wire dma_write_addr3_to_bank6      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr3_to_bank6       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank6   =  dma_write_addr3_to_bank6  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank6    =  write_request3_to_bank6   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank6    =  dma_read_addr3_to_bank6   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank6     =  read_request3_to_bank6    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank7
  wire dma_write_addr3_to_bank7      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr3_to_bank7       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank7   =  dma_write_addr3_to_bank7  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank7    =  write_request3_to_bank7   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank7    =  dma_read_addr3_to_bank7   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank7     =  read_request3_to_bank7    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank8
  wire dma_write_addr3_to_bank8      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr3_to_bank8       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank8   =  dma_write_addr3_to_bank8  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank8    =  write_request3_to_bank8   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank8    =  dma_read_addr3_to_bank8   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank8     =  read_request3_to_bank8    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank9
  wire dma_write_addr3_to_bank9      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr3_to_bank9       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank9   =  dma_write_addr3_to_bank9  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank9    =  write_request3_to_bank9   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank9    =  dma_read_addr3_to_bank9   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank9     =  read_request3_to_bank9    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank10
  wire dma_write_addr3_to_bank10      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr3_to_bank10       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank10   =  dma_write_addr3_to_bank10  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank10    =  write_request3_to_bank10   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank10    =  dma_read_addr3_to_bank10   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank10     =  read_request3_to_bank10    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank11
  wire dma_write_addr3_to_bank11      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr3_to_bank11       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank11   =  dma_write_addr3_to_bank11  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank11    =  write_request3_to_bank11   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank11    =  dma_read_addr3_to_bank11   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank11     =  read_request3_to_bank11    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank12
  wire dma_write_addr3_to_bank12      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr3_to_bank12       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank12   =  dma_write_addr3_to_bank12  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank12    =  write_request3_to_bank12   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank12    =  dma_read_addr3_to_bank12   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank12     =  read_request3_to_bank12    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank13
  wire dma_write_addr3_to_bank13      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr3_to_bank13       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank13   =  dma_write_addr3_to_bank13  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank13    =  write_request3_to_bank13   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank13    =  dma_read_addr3_to_bank13   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank13     =  read_request3_to_bank13    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank14
  wire dma_write_addr3_to_bank14      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr3_to_bank14       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank14   =  dma_write_addr3_to_bank14  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank14    =  write_request3_to_bank14   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank14    =  dma_read_addr3_to_bank14   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank14     =  read_request3_to_bank14    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank15
  wire dma_write_addr3_to_bank15      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr3_to_bank15       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank15   =  dma_write_addr3_to_bank15  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank15    =  write_request3_to_bank15   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank15    =  dma_read_addr3_to_bank15   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank15     =  read_request3_to_bank15    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank16
  wire dma_write_addr3_to_bank16      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr3_to_bank16       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank16   =  dma_write_addr3_to_bank16  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank16    =  write_request3_to_bank16   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank16    =  dma_read_addr3_to_bank16   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank16     =  read_request3_to_bank16    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank17
  wire dma_write_addr3_to_bank17      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr3_to_bank17       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank17   =  dma_write_addr3_to_bank17  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank17    =  write_request3_to_bank17   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank17    =  dma_read_addr3_to_bank17   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank17     =  read_request3_to_bank17    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank18
  wire dma_write_addr3_to_bank18      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr3_to_bank18       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank18   =  dma_write_addr3_to_bank18  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank18    =  write_request3_to_bank18   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank18    =  dma_read_addr3_to_bank18   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank18     =  read_request3_to_bank18    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank19
  wire dma_write_addr3_to_bank19      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr3_to_bank19       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank19   =  dma_write_addr3_to_bank19  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank19    =  write_request3_to_bank19   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank19    =  dma_read_addr3_to_bank19   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank19     =  read_request3_to_bank19    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank20
  wire dma_write_addr3_to_bank20      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr3_to_bank20       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank20   =  dma_write_addr3_to_bank20  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank20    =  write_request3_to_bank20   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank20    =  dma_read_addr3_to_bank20   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank20     =  read_request3_to_bank20    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank21
  wire dma_write_addr3_to_bank21      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr3_to_bank21       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank21   =  dma_write_addr3_to_bank21  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank21    =  write_request3_to_bank21   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank21    =  dma_read_addr3_to_bank21   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank21     =  read_request3_to_bank21    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank22
  wire dma_write_addr3_to_bank22      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr3_to_bank22       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank22   =  dma_write_addr3_to_bank22  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank22    =  write_request3_to_bank22   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank22    =  dma_read_addr3_to_bank22   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank22     =  read_request3_to_bank22    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank23
  wire dma_write_addr3_to_bank23      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr3_to_bank23       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank23   =  dma_write_addr3_to_bank23  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank23    =  write_request3_to_bank23   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank23    =  dma_read_addr3_to_bank23   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank23     =  read_request3_to_bank23    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank24
  wire dma_write_addr3_to_bank24      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr3_to_bank24       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank24   =  dma_write_addr3_to_bank24  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank24    =  write_request3_to_bank24   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank24    =  dma_read_addr3_to_bank24   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank24     =  read_request3_to_bank24    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank25
  wire dma_write_addr3_to_bank25      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr3_to_bank25       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank25   =  dma_write_addr3_to_bank25  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank25    =  write_request3_to_bank25   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank25    =  dma_read_addr3_to_bank25   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank25     =  read_request3_to_bank25    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank26
  wire dma_write_addr3_to_bank26      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr3_to_bank26       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank26   =  dma_write_addr3_to_bank26  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank26    =  write_request3_to_bank26   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank26    =  dma_read_addr3_to_bank26   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank26     =  read_request3_to_bank26    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank27
  wire dma_write_addr3_to_bank27      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr3_to_bank27       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank27   =  dma_write_addr3_to_bank27  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank27    =  write_request3_to_bank27   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank27    =  dma_read_addr3_to_bank27   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank27     =  read_request3_to_bank27    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank28
  wire dma_write_addr3_to_bank28      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr3_to_bank28       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank28   =  dma_write_addr3_to_bank28  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank28    =  write_request3_to_bank28   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank28    =  dma_read_addr3_to_bank28   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank28     =  read_request3_to_bank28    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank29
  wire dma_write_addr3_to_bank29      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr3_to_bank29       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank29   =  dma_write_addr3_to_bank29  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank29    =  write_request3_to_bank29   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank29    =  dma_read_addr3_to_bank29   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank29     =  read_request3_to_bank29    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank30
  wire dma_write_addr3_to_bank30      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr3_to_bank30       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank30   =  dma_write_addr3_to_bank30  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank30    =  write_request3_to_bank30   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank30    =  dma_read_addr3_to_bank30   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank30     =  read_request3_to_bank30    & memc__dma__read_ready3   ;                                         
  // DMA 3, bank31
  wire dma_write_addr3_to_bank31      =  (dma__memc__write_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr3_to_bank31       =  (dma__memc__read_address3[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank31   =  dma_write_addr3_to_bank31  & dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank31    =  write_request3_to_bank31   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank31    =  dma_read_addr3_to_bank31   & dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank31     =  read_request3_to_bank31    & memc__dma__read_ready3   ;                                         
  // DMA 4
  wire read_pause4     =  dma__memc__read_pause4   ;  
  // DMA 4, bank0
  wire dma_write_addr4_to_bank0      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr4_to_bank0       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank0   =  dma_write_addr4_to_bank0  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank0    =  write_request4_to_bank0   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank0    =  dma_read_addr4_to_bank0   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank0     =  read_request4_to_bank0    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank1
  wire dma_write_addr4_to_bank1      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr4_to_bank1       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank1   =  dma_write_addr4_to_bank1  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank1    =  write_request4_to_bank1   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank1    =  dma_read_addr4_to_bank1   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank1     =  read_request4_to_bank1    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank2
  wire dma_write_addr4_to_bank2      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr4_to_bank2       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank2   =  dma_write_addr4_to_bank2  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank2    =  write_request4_to_bank2   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank2    =  dma_read_addr4_to_bank2   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank2     =  read_request4_to_bank2    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank3
  wire dma_write_addr4_to_bank3      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr4_to_bank3       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank3   =  dma_write_addr4_to_bank3  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank3    =  write_request4_to_bank3   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank3    =  dma_read_addr4_to_bank3   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank3     =  read_request4_to_bank3    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank4
  wire dma_write_addr4_to_bank4      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr4_to_bank4       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank4   =  dma_write_addr4_to_bank4  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank4    =  write_request4_to_bank4   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank4    =  dma_read_addr4_to_bank4   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank4     =  read_request4_to_bank4    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank5
  wire dma_write_addr4_to_bank5      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr4_to_bank5       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank5   =  dma_write_addr4_to_bank5  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank5    =  write_request4_to_bank5   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank5    =  dma_read_addr4_to_bank5   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank5     =  read_request4_to_bank5    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank6
  wire dma_write_addr4_to_bank6      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr4_to_bank6       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank6   =  dma_write_addr4_to_bank6  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank6    =  write_request4_to_bank6   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank6    =  dma_read_addr4_to_bank6   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank6     =  read_request4_to_bank6    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank7
  wire dma_write_addr4_to_bank7      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr4_to_bank7       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank7   =  dma_write_addr4_to_bank7  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank7    =  write_request4_to_bank7   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank7    =  dma_read_addr4_to_bank7   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank7     =  read_request4_to_bank7    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank8
  wire dma_write_addr4_to_bank8      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr4_to_bank8       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank8   =  dma_write_addr4_to_bank8  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank8    =  write_request4_to_bank8   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank8    =  dma_read_addr4_to_bank8   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank8     =  read_request4_to_bank8    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank9
  wire dma_write_addr4_to_bank9      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr4_to_bank9       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank9   =  dma_write_addr4_to_bank9  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank9    =  write_request4_to_bank9   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank9    =  dma_read_addr4_to_bank9   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank9     =  read_request4_to_bank9    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank10
  wire dma_write_addr4_to_bank10      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr4_to_bank10       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank10   =  dma_write_addr4_to_bank10  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank10    =  write_request4_to_bank10   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank10    =  dma_read_addr4_to_bank10   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank10     =  read_request4_to_bank10    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank11
  wire dma_write_addr4_to_bank11      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr4_to_bank11       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank11   =  dma_write_addr4_to_bank11  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank11    =  write_request4_to_bank11   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank11    =  dma_read_addr4_to_bank11   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank11     =  read_request4_to_bank11    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank12
  wire dma_write_addr4_to_bank12      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr4_to_bank12       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank12   =  dma_write_addr4_to_bank12  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank12    =  write_request4_to_bank12   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank12    =  dma_read_addr4_to_bank12   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank12     =  read_request4_to_bank12    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank13
  wire dma_write_addr4_to_bank13      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr4_to_bank13       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank13   =  dma_write_addr4_to_bank13  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank13    =  write_request4_to_bank13   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank13    =  dma_read_addr4_to_bank13   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank13     =  read_request4_to_bank13    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank14
  wire dma_write_addr4_to_bank14      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr4_to_bank14       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank14   =  dma_write_addr4_to_bank14  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank14    =  write_request4_to_bank14   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank14    =  dma_read_addr4_to_bank14   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank14     =  read_request4_to_bank14    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank15
  wire dma_write_addr4_to_bank15      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr4_to_bank15       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank15   =  dma_write_addr4_to_bank15  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank15    =  write_request4_to_bank15   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank15    =  dma_read_addr4_to_bank15   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank15     =  read_request4_to_bank15    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank16
  wire dma_write_addr4_to_bank16      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr4_to_bank16       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank16   =  dma_write_addr4_to_bank16  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank16    =  write_request4_to_bank16   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank16    =  dma_read_addr4_to_bank16   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank16     =  read_request4_to_bank16    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank17
  wire dma_write_addr4_to_bank17      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr4_to_bank17       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank17   =  dma_write_addr4_to_bank17  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank17    =  write_request4_to_bank17   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank17    =  dma_read_addr4_to_bank17   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank17     =  read_request4_to_bank17    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank18
  wire dma_write_addr4_to_bank18      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr4_to_bank18       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank18   =  dma_write_addr4_to_bank18  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank18    =  write_request4_to_bank18   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank18    =  dma_read_addr4_to_bank18   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank18     =  read_request4_to_bank18    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank19
  wire dma_write_addr4_to_bank19      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr4_to_bank19       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank19   =  dma_write_addr4_to_bank19  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank19    =  write_request4_to_bank19   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank19    =  dma_read_addr4_to_bank19   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank19     =  read_request4_to_bank19    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank20
  wire dma_write_addr4_to_bank20      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr4_to_bank20       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank20   =  dma_write_addr4_to_bank20  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank20    =  write_request4_to_bank20   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank20    =  dma_read_addr4_to_bank20   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank20     =  read_request4_to_bank20    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank21
  wire dma_write_addr4_to_bank21      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr4_to_bank21       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank21   =  dma_write_addr4_to_bank21  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank21    =  write_request4_to_bank21   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank21    =  dma_read_addr4_to_bank21   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank21     =  read_request4_to_bank21    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank22
  wire dma_write_addr4_to_bank22      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr4_to_bank22       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank22   =  dma_write_addr4_to_bank22  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank22    =  write_request4_to_bank22   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank22    =  dma_read_addr4_to_bank22   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank22     =  read_request4_to_bank22    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank23
  wire dma_write_addr4_to_bank23      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr4_to_bank23       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank23   =  dma_write_addr4_to_bank23  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank23    =  write_request4_to_bank23   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank23    =  dma_read_addr4_to_bank23   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank23     =  read_request4_to_bank23    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank24
  wire dma_write_addr4_to_bank24      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr4_to_bank24       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank24   =  dma_write_addr4_to_bank24  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank24    =  write_request4_to_bank24   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank24    =  dma_read_addr4_to_bank24   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank24     =  read_request4_to_bank24    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank25
  wire dma_write_addr4_to_bank25      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr4_to_bank25       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank25   =  dma_write_addr4_to_bank25  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank25    =  write_request4_to_bank25   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank25    =  dma_read_addr4_to_bank25   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank25     =  read_request4_to_bank25    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank26
  wire dma_write_addr4_to_bank26      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr4_to_bank26       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank26   =  dma_write_addr4_to_bank26  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank26    =  write_request4_to_bank26   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank26    =  dma_read_addr4_to_bank26   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank26     =  read_request4_to_bank26    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank27
  wire dma_write_addr4_to_bank27      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr4_to_bank27       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank27   =  dma_write_addr4_to_bank27  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank27    =  write_request4_to_bank27   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank27    =  dma_read_addr4_to_bank27   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank27     =  read_request4_to_bank27    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank28
  wire dma_write_addr4_to_bank28      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr4_to_bank28       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank28   =  dma_write_addr4_to_bank28  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank28    =  write_request4_to_bank28   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank28    =  dma_read_addr4_to_bank28   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank28     =  read_request4_to_bank28    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank29
  wire dma_write_addr4_to_bank29      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr4_to_bank29       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank29   =  dma_write_addr4_to_bank29  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank29    =  write_request4_to_bank29   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank29    =  dma_read_addr4_to_bank29   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank29     =  read_request4_to_bank29    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank30
  wire dma_write_addr4_to_bank30      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr4_to_bank30       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank30   =  dma_write_addr4_to_bank30  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank30    =  write_request4_to_bank30   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank30    =  dma_read_addr4_to_bank30   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank30     =  read_request4_to_bank30    & memc__dma__read_ready4   ;                                         
  // DMA 4, bank31
  wire dma_write_addr4_to_bank31      =  (dma__memc__write_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr4_to_bank31       =  (dma__memc__read_address4[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank31   =  dma_write_addr4_to_bank31  & dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank31    =  write_request4_to_bank31   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank31    =  dma_read_addr4_to_bank31   & dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank31     =  read_request4_to_bank31    & memc__dma__read_ready4   ;                                         
  // DMA 5
  wire read_pause5     =  dma__memc__read_pause5   ;  
  // DMA 5, bank0
  wire dma_write_addr5_to_bank0      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr5_to_bank0       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank0   =  dma_write_addr5_to_bank0  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank0    =  write_request5_to_bank0   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank0    =  dma_read_addr5_to_bank0   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank0     =  read_request5_to_bank0    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank1
  wire dma_write_addr5_to_bank1      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr5_to_bank1       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank1   =  dma_write_addr5_to_bank1  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank1    =  write_request5_to_bank1   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank1    =  dma_read_addr5_to_bank1   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank1     =  read_request5_to_bank1    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank2
  wire dma_write_addr5_to_bank2      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr5_to_bank2       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank2   =  dma_write_addr5_to_bank2  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank2    =  write_request5_to_bank2   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank2    =  dma_read_addr5_to_bank2   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank2     =  read_request5_to_bank2    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank3
  wire dma_write_addr5_to_bank3      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr5_to_bank3       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank3   =  dma_write_addr5_to_bank3  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank3    =  write_request5_to_bank3   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank3    =  dma_read_addr5_to_bank3   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank3     =  read_request5_to_bank3    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank4
  wire dma_write_addr5_to_bank4      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr5_to_bank4       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank4   =  dma_write_addr5_to_bank4  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank4    =  write_request5_to_bank4   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank4    =  dma_read_addr5_to_bank4   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank4     =  read_request5_to_bank4    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank5
  wire dma_write_addr5_to_bank5      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr5_to_bank5       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank5   =  dma_write_addr5_to_bank5  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank5    =  write_request5_to_bank5   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank5    =  dma_read_addr5_to_bank5   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank5     =  read_request5_to_bank5    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank6
  wire dma_write_addr5_to_bank6      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr5_to_bank6       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank6   =  dma_write_addr5_to_bank6  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank6    =  write_request5_to_bank6   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank6    =  dma_read_addr5_to_bank6   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank6     =  read_request5_to_bank6    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank7
  wire dma_write_addr5_to_bank7      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr5_to_bank7       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank7   =  dma_write_addr5_to_bank7  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank7    =  write_request5_to_bank7   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank7    =  dma_read_addr5_to_bank7   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank7     =  read_request5_to_bank7    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank8
  wire dma_write_addr5_to_bank8      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr5_to_bank8       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank8   =  dma_write_addr5_to_bank8  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank8    =  write_request5_to_bank8   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank8    =  dma_read_addr5_to_bank8   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank8     =  read_request5_to_bank8    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank9
  wire dma_write_addr5_to_bank9      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr5_to_bank9       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank9   =  dma_write_addr5_to_bank9  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank9    =  write_request5_to_bank9   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank9    =  dma_read_addr5_to_bank9   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank9     =  read_request5_to_bank9    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank10
  wire dma_write_addr5_to_bank10      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr5_to_bank10       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank10   =  dma_write_addr5_to_bank10  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank10    =  write_request5_to_bank10   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank10    =  dma_read_addr5_to_bank10   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank10     =  read_request5_to_bank10    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank11
  wire dma_write_addr5_to_bank11      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr5_to_bank11       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank11   =  dma_write_addr5_to_bank11  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank11    =  write_request5_to_bank11   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank11    =  dma_read_addr5_to_bank11   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank11     =  read_request5_to_bank11    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank12
  wire dma_write_addr5_to_bank12      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr5_to_bank12       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank12   =  dma_write_addr5_to_bank12  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank12    =  write_request5_to_bank12   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank12    =  dma_read_addr5_to_bank12   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank12     =  read_request5_to_bank12    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank13
  wire dma_write_addr5_to_bank13      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr5_to_bank13       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank13   =  dma_write_addr5_to_bank13  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank13    =  write_request5_to_bank13   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank13    =  dma_read_addr5_to_bank13   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank13     =  read_request5_to_bank13    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank14
  wire dma_write_addr5_to_bank14      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr5_to_bank14       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank14   =  dma_write_addr5_to_bank14  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank14    =  write_request5_to_bank14   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank14    =  dma_read_addr5_to_bank14   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank14     =  read_request5_to_bank14    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank15
  wire dma_write_addr5_to_bank15      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr5_to_bank15       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank15   =  dma_write_addr5_to_bank15  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank15    =  write_request5_to_bank15   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank15    =  dma_read_addr5_to_bank15   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank15     =  read_request5_to_bank15    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank16
  wire dma_write_addr5_to_bank16      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr5_to_bank16       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank16   =  dma_write_addr5_to_bank16  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank16    =  write_request5_to_bank16   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank16    =  dma_read_addr5_to_bank16   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank16     =  read_request5_to_bank16    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank17
  wire dma_write_addr5_to_bank17      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr5_to_bank17       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank17   =  dma_write_addr5_to_bank17  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank17    =  write_request5_to_bank17   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank17    =  dma_read_addr5_to_bank17   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank17     =  read_request5_to_bank17    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank18
  wire dma_write_addr5_to_bank18      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr5_to_bank18       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank18   =  dma_write_addr5_to_bank18  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank18    =  write_request5_to_bank18   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank18    =  dma_read_addr5_to_bank18   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank18     =  read_request5_to_bank18    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank19
  wire dma_write_addr5_to_bank19      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr5_to_bank19       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank19   =  dma_write_addr5_to_bank19  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank19    =  write_request5_to_bank19   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank19    =  dma_read_addr5_to_bank19   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank19     =  read_request5_to_bank19    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank20
  wire dma_write_addr5_to_bank20      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr5_to_bank20       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank20   =  dma_write_addr5_to_bank20  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank20    =  write_request5_to_bank20   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank20    =  dma_read_addr5_to_bank20   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank20     =  read_request5_to_bank20    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank21
  wire dma_write_addr5_to_bank21      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr5_to_bank21       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank21   =  dma_write_addr5_to_bank21  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank21    =  write_request5_to_bank21   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank21    =  dma_read_addr5_to_bank21   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank21     =  read_request5_to_bank21    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank22
  wire dma_write_addr5_to_bank22      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr5_to_bank22       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank22   =  dma_write_addr5_to_bank22  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank22    =  write_request5_to_bank22   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank22    =  dma_read_addr5_to_bank22   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank22     =  read_request5_to_bank22    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank23
  wire dma_write_addr5_to_bank23      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr5_to_bank23       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank23   =  dma_write_addr5_to_bank23  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank23    =  write_request5_to_bank23   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank23    =  dma_read_addr5_to_bank23   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank23     =  read_request5_to_bank23    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank24
  wire dma_write_addr5_to_bank24      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr5_to_bank24       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank24   =  dma_write_addr5_to_bank24  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank24    =  write_request5_to_bank24   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank24    =  dma_read_addr5_to_bank24   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank24     =  read_request5_to_bank24    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank25
  wire dma_write_addr5_to_bank25      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr5_to_bank25       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank25   =  dma_write_addr5_to_bank25  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank25    =  write_request5_to_bank25   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank25    =  dma_read_addr5_to_bank25   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank25     =  read_request5_to_bank25    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank26
  wire dma_write_addr5_to_bank26      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr5_to_bank26       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank26   =  dma_write_addr5_to_bank26  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank26    =  write_request5_to_bank26   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank26    =  dma_read_addr5_to_bank26   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank26     =  read_request5_to_bank26    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank27
  wire dma_write_addr5_to_bank27      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr5_to_bank27       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank27   =  dma_write_addr5_to_bank27  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank27    =  write_request5_to_bank27   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank27    =  dma_read_addr5_to_bank27   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank27     =  read_request5_to_bank27    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank28
  wire dma_write_addr5_to_bank28      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr5_to_bank28       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank28   =  dma_write_addr5_to_bank28  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank28    =  write_request5_to_bank28   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank28    =  dma_read_addr5_to_bank28   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank28     =  read_request5_to_bank28    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank29
  wire dma_write_addr5_to_bank29      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr5_to_bank29       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank29   =  dma_write_addr5_to_bank29  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank29    =  write_request5_to_bank29   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank29    =  dma_read_addr5_to_bank29   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank29     =  read_request5_to_bank29    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank30
  wire dma_write_addr5_to_bank30      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr5_to_bank30       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank30   =  dma_write_addr5_to_bank30  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank30    =  write_request5_to_bank30   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank30    =  dma_read_addr5_to_bank30   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank30     =  read_request5_to_bank30    & memc__dma__read_ready5   ;                                         
  // DMA 5, bank31
  wire dma_write_addr5_to_bank31      =  (dma__memc__write_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr5_to_bank31       =  (dma__memc__read_address5[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank31   =  dma_write_addr5_to_bank31  & dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank31    =  write_request5_to_bank31   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank31    =  dma_read_addr5_to_bank31   & dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank31     =  read_request5_to_bank31    & memc__dma__read_ready5   ;                                         
  // DMA 6
  wire read_pause6     =  dma__memc__read_pause6   ;  
  // DMA 6, bank0
  wire dma_write_addr6_to_bank0      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr6_to_bank0       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank0   =  dma_write_addr6_to_bank0  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank0    =  write_request6_to_bank0   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank0    =  dma_read_addr6_to_bank0   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank0     =  read_request6_to_bank0    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank1
  wire dma_write_addr6_to_bank1      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr6_to_bank1       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank1   =  dma_write_addr6_to_bank1  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank1    =  write_request6_to_bank1   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank1    =  dma_read_addr6_to_bank1   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank1     =  read_request6_to_bank1    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank2
  wire dma_write_addr6_to_bank2      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr6_to_bank2       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank2   =  dma_write_addr6_to_bank2  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank2    =  write_request6_to_bank2   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank2    =  dma_read_addr6_to_bank2   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank2     =  read_request6_to_bank2    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank3
  wire dma_write_addr6_to_bank3      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr6_to_bank3       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank3   =  dma_write_addr6_to_bank3  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank3    =  write_request6_to_bank3   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank3    =  dma_read_addr6_to_bank3   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank3     =  read_request6_to_bank3    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank4
  wire dma_write_addr6_to_bank4      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr6_to_bank4       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank4   =  dma_write_addr6_to_bank4  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank4    =  write_request6_to_bank4   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank4    =  dma_read_addr6_to_bank4   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank4     =  read_request6_to_bank4    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank5
  wire dma_write_addr6_to_bank5      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr6_to_bank5       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank5   =  dma_write_addr6_to_bank5  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank5    =  write_request6_to_bank5   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank5    =  dma_read_addr6_to_bank5   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank5     =  read_request6_to_bank5    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank6
  wire dma_write_addr6_to_bank6      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr6_to_bank6       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank6   =  dma_write_addr6_to_bank6  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank6    =  write_request6_to_bank6   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank6    =  dma_read_addr6_to_bank6   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank6     =  read_request6_to_bank6    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank7
  wire dma_write_addr6_to_bank7      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr6_to_bank7       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank7   =  dma_write_addr6_to_bank7  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank7    =  write_request6_to_bank7   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank7    =  dma_read_addr6_to_bank7   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank7     =  read_request6_to_bank7    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank8
  wire dma_write_addr6_to_bank8      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr6_to_bank8       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank8   =  dma_write_addr6_to_bank8  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank8    =  write_request6_to_bank8   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank8    =  dma_read_addr6_to_bank8   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank8     =  read_request6_to_bank8    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank9
  wire dma_write_addr6_to_bank9      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr6_to_bank9       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank9   =  dma_write_addr6_to_bank9  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank9    =  write_request6_to_bank9   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank9    =  dma_read_addr6_to_bank9   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank9     =  read_request6_to_bank9    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank10
  wire dma_write_addr6_to_bank10      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr6_to_bank10       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank10   =  dma_write_addr6_to_bank10  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank10    =  write_request6_to_bank10   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank10    =  dma_read_addr6_to_bank10   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank10     =  read_request6_to_bank10    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank11
  wire dma_write_addr6_to_bank11      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr6_to_bank11       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank11   =  dma_write_addr6_to_bank11  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank11    =  write_request6_to_bank11   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank11    =  dma_read_addr6_to_bank11   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank11     =  read_request6_to_bank11    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank12
  wire dma_write_addr6_to_bank12      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr6_to_bank12       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank12   =  dma_write_addr6_to_bank12  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank12    =  write_request6_to_bank12   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank12    =  dma_read_addr6_to_bank12   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank12     =  read_request6_to_bank12    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank13
  wire dma_write_addr6_to_bank13      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr6_to_bank13       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank13   =  dma_write_addr6_to_bank13  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank13    =  write_request6_to_bank13   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank13    =  dma_read_addr6_to_bank13   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank13     =  read_request6_to_bank13    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank14
  wire dma_write_addr6_to_bank14      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr6_to_bank14       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank14   =  dma_write_addr6_to_bank14  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank14    =  write_request6_to_bank14   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank14    =  dma_read_addr6_to_bank14   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank14     =  read_request6_to_bank14    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank15
  wire dma_write_addr6_to_bank15      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr6_to_bank15       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank15   =  dma_write_addr6_to_bank15  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank15    =  write_request6_to_bank15   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank15    =  dma_read_addr6_to_bank15   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank15     =  read_request6_to_bank15    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank16
  wire dma_write_addr6_to_bank16      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr6_to_bank16       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank16   =  dma_write_addr6_to_bank16  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank16    =  write_request6_to_bank16   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank16    =  dma_read_addr6_to_bank16   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank16     =  read_request6_to_bank16    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank17
  wire dma_write_addr6_to_bank17      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr6_to_bank17       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank17   =  dma_write_addr6_to_bank17  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank17    =  write_request6_to_bank17   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank17    =  dma_read_addr6_to_bank17   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank17     =  read_request6_to_bank17    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank18
  wire dma_write_addr6_to_bank18      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr6_to_bank18       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank18   =  dma_write_addr6_to_bank18  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank18    =  write_request6_to_bank18   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank18    =  dma_read_addr6_to_bank18   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank18     =  read_request6_to_bank18    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank19
  wire dma_write_addr6_to_bank19      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr6_to_bank19       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank19   =  dma_write_addr6_to_bank19  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank19    =  write_request6_to_bank19   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank19    =  dma_read_addr6_to_bank19   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank19     =  read_request6_to_bank19    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank20
  wire dma_write_addr6_to_bank20      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr6_to_bank20       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank20   =  dma_write_addr6_to_bank20  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank20    =  write_request6_to_bank20   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank20    =  dma_read_addr6_to_bank20   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank20     =  read_request6_to_bank20    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank21
  wire dma_write_addr6_to_bank21      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr6_to_bank21       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank21   =  dma_write_addr6_to_bank21  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank21    =  write_request6_to_bank21   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank21    =  dma_read_addr6_to_bank21   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank21     =  read_request6_to_bank21    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank22
  wire dma_write_addr6_to_bank22      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr6_to_bank22       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank22   =  dma_write_addr6_to_bank22  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank22    =  write_request6_to_bank22   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank22    =  dma_read_addr6_to_bank22   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank22     =  read_request6_to_bank22    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank23
  wire dma_write_addr6_to_bank23      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr6_to_bank23       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank23   =  dma_write_addr6_to_bank23  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank23    =  write_request6_to_bank23   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank23    =  dma_read_addr6_to_bank23   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank23     =  read_request6_to_bank23    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank24
  wire dma_write_addr6_to_bank24      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr6_to_bank24       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank24   =  dma_write_addr6_to_bank24  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank24    =  write_request6_to_bank24   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank24    =  dma_read_addr6_to_bank24   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank24     =  read_request6_to_bank24    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank25
  wire dma_write_addr6_to_bank25      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr6_to_bank25       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank25   =  dma_write_addr6_to_bank25  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank25    =  write_request6_to_bank25   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank25    =  dma_read_addr6_to_bank25   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank25     =  read_request6_to_bank25    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank26
  wire dma_write_addr6_to_bank26      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr6_to_bank26       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank26   =  dma_write_addr6_to_bank26  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank26    =  write_request6_to_bank26   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank26    =  dma_read_addr6_to_bank26   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank26     =  read_request6_to_bank26    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank27
  wire dma_write_addr6_to_bank27      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr6_to_bank27       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank27   =  dma_write_addr6_to_bank27  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank27    =  write_request6_to_bank27   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank27    =  dma_read_addr6_to_bank27   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank27     =  read_request6_to_bank27    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank28
  wire dma_write_addr6_to_bank28      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr6_to_bank28       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank28   =  dma_write_addr6_to_bank28  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank28    =  write_request6_to_bank28   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank28    =  dma_read_addr6_to_bank28   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank28     =  read_request6_to_bank28    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank29
  wire dma_write_addr6_to_bank29      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr6_to_bank29       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank29   =  dma_write_addr6_to_bank29  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank29    =  write_request6_to_bank29   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank29    =  dma_read_addr6_to_bank29   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank29     =  read_request6_to_bank29    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank30
  wire dma_write_addr6_to_bank30      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr6_to_bank30       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank30   =  dma_write_addr6_to_bank30  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank30    =  write_request6_to_bank30   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank30    =  dma_read_addr6_to_bank30   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank30     =  read_request6_to_bank30    & memc__dma__read_ready6   ;                                         
  // DMA 6, bank31
  wire dma_write_addr6_to_bank31      =  (dma__memc__write_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr6_to_bank31       =  (dma__memc__read_address6[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank31   =  dma_write_addr6_to_bank31  & dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank31    =  write_request6_to_bank31   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank31    =  dma_read_addr6_to_bank31   & dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank31     =  read_request6_to_bank31    & memc__dma__read_ready6   ;                                         
  // DMA 7
  wire read_pause7     =  dma__memc__read_pause7   ;  
  // DMA 7, bank0
  wire dma_write_addr7_to_bank0      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr7_to_bank0       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank0   =  dma_write_addr7_to_bank0  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank0    =  write_request7_to_bank0   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank0    =  dma_read_addr7_to_bank0   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank0     =  read_request7_to_bank0    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank1
  wire dma_write_addr7_to_bank1      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr7_to_bank1       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank1   =  dma_write_addr7_to_bank1  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank1    =  write_request7_to_bank1   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank1    =  dma_read_addr7_to_bank1   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank1     =  read_request7_to_bank1    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank2
  wire dma_write_addr7_to_bank2      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr7_to_bank2       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank2   =  dma_write_addr7_to_bank2  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank2    =  write_request7_to_bank2   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank2    =  dma_read_addr7_to_bank2   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank2     =  read_request7_to_bank2    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank3
  wire dma_write_addr7_to_bank3      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr7_to_bank3       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank3   =  dma_write_addr7_to_bank3  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank3    =  write_request7_to_bank3   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank3    =  dma_read_addr7_to_bank3   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank3     =  read_request7_to_bank3    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank4
  wire dma_write_addr7_to_bank4      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr7_to_bank4       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank4   =  dma_write_addr7_to_bank4  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank4    =  write_request7_to_bank4   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank4    =  dma_read_addr7_to_bank4   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank4     =  read_request7_to_bank4    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank5
  wire dma_write_addr7_to_bank5      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr7_to_bank5       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank5   =  dma_write_addr7_to_bank5  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank5    =  write_request7_to_bank5   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank5    =  dma_read_addr7_to_bank5   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank5     =  read_request7_to_bank5    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank6
  wire dma_write_addr7_to_bank6      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr7_to_bank6       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank6   =  dma_write_addr7_to_bank6  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank6    =  write_request7_to_bank6   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank6    =  dma_read_addr7_to_bank6   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank6     =  read_request7_to_bank6    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank7
  wire dma_write_addr7_to_bank7      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr7_to_bank7       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank7   =  dma_write_addr7_to_bank7  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank7    =  write_request7_to_bank7   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank7    =  dma_read_addr7_to_bank7   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank7     =  read_request7_to_bank7    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank8
  wire dma_write_addr7_to_bank8      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr7_to_bank8       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank8   =  dma_write_addr7_to_bank8  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank8    =  write_request7_to_bank8   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank8    =  dma_read_addr7_to_bank8   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank8     =  read_request7_to_bank8    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank9
  wire dma_write_addr7_to_bank9      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr7_to_bank9       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank9   =  dma_write_addr7_to_bank9  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank9    =  write_request7_to_bank9   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank9    =  dma_read_addr7_to_bank9   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank9     =  read_request7_to_bank9    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank10
  wire dma_write_addr7_to_bank10      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr7_to_bank10       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank10   =  dma_write_addr7_to_bank10  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank10    =  write_request7_to_bank10   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank10    =  dma_read_addr7_to_bank10   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank10     =  read_request7_to_bank10    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank11
  wire dma_write_addr7_to_bank11      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr7_to_bank11       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank11   =  dma_write_addr7_to_bank11  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank11    =  write_request7_to_bank11   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank11    =  dma_read_addr7_to_bank11   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank11     =  read_request7_to_bank11    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank12
  wire dma_write_addr7_to_bank12      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr7_to_bank12       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank12   =  dma_write_addr7_to_bank12  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank12    =  write_request7_to_bank12   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank12    =  dma_read_addr7_to_bank12   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank12     =  read_request7_to_bank12    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank13
  wire dma_write_addr7_to_bank13      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr7_to_bank13       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank13   =  dma_write_addr7_to_bank13  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank13    =  write_request7_to_bank13   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank13    =  dma_read_addr7_to_bank13   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank13     =  read_request7_to_bank13    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank14
  wire dma_write_addr7_to_bank14      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr7_to_bank14       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank14   =  dma_write_addr7_to_bank14  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank14    =  write_request7_to_bank14   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank14    =  dma_read_addr7_to_bank14   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank14     =  read_request7_to_bank14    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank15
  wire dma_write_addr7_to_bank15      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr7_to_bank15       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank15   =  dma_write_addr7_to_bank15  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank15    =  write_request7_to_bank15   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank15    =  dma_read_addr7_to_bank15   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank15     =  read_request7_to_bank15    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank16
  wire dma_write_addr7_to_bank16      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr7_to_bank16       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank16   =  dma_write_addr7_to_bank16  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank16    =  write_request7_to_bank16   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank16    =  dma_read_addr7_to_bank16   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank16     =  read_request7_to_bank16    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank17
  wire dma_write_addr7_to_bank17      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr7_to_bank17       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank17   =  dma_write_addr7_to_bank17  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank17    =  write_request7_to_bank17   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank17    =  dma_read_addr7_to_bank17   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank17     =  read_request7_to_bank17    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank18
  wire dma_write_addr7_to_bank18      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr7_to_bank18       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank18   =  dma_write_addr7_to_bank18  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank18    =  write_request7_to_bank18   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank18    =  dma_read_addr7_to_bank18   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank18     =  read_request7_to_bank18    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank19
  wire dma_write_addr7_to_bank19      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr7_to_bank19       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank19   =  dma_write_addr7_to_bank19  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank19    =  write_request7_to_bank19   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank19    =  dma_read_addr7_to_bank19   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank19     =  read_request7_to_bank19    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank20
  wire dma_write_addr7_to_bank20      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr7_to_bank20       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank20   =  dma_write_addr7_to_bank20  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank20    =  write_request7_to_bank20   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank20    =  dma_read_addr7_to_bank20   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank20     =  read_request7_to_bank20    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank21
  wire dma_write_addr7_to_bank21      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr7_to_bank21       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank21   =  dma_write_addr7_to_bank21  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank21    =  write_request7_to_bank21   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank21    =  dma_read_addr7_to_bank21   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank21     =  read_request7_to_bank21    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank22
  wire dma_write_addr7_to_bank22      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr7_to_bank22       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank22   =  dma_write_addr7_to_bank22  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank22    =  write_request7_to_bank22   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank22    =  dma_read_addr7_to_bank22   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank22     =  read_request7_to_bank22    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank23
  wire dma_write_addr7_to_bank23      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr7_to_bank23       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank23   =  dma_write_addr7_to_bank23  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank23    =  write_request7_to_bank23   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank23    =  dma_read_addr7_to_bank23   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank23     =  read_request7_to_bank23    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank24
  wire dma_write_addr7_to_bank24      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr7_to_bank24       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank24   =  dma_write_addr7_to_bank24  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank24    =  write_request7_to_bank24   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank24    =  dma_read_addr7_to_bank24   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank24     =  read_request7_to_bank24    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank25
  wire dma_write_addr7_to_bank25      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr7_to_bank25       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank25   =  dma_write_addr7_to_bank25  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank25    =  write_request7_to_bank25   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank25    =  dma_read_addr7_to_bank25   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank25     =  read_request7_to_bank25    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank26
  wire dma_write_addr7_to_bank26      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr7_to_bank26       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank26   =  dma_write_addr7_to_bank26  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank26    =  write_request7_to_bank26   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank26    =  dma_read_addr7_to_bank26   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank26     =  read_request7_to_bank26    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank27
  wire dma_write_addr7_to_bank27      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr7_to_bank27       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank27   =  dma_write_addr7_to_bank27  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank27    =  write_request7_to_bank27   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank27    =  dma_read_addr7_to_bank27   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank27     =  read_request7_to_bank27    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank28
  wire dma_write_addr7_to_bank28      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr7_to_bank28       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank28   =  dma_write_addr7_to_bank28  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank28    =  write_request7_to_bank28   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank28    =  dma_read_addr7_to_bank28   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank28     =  read_request7_to_bank28    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank29
  wire dma_write_addr7_to_bank29      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr7_to_bank29       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank29   =  dma_write_addr7_to_bank29  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank29    =  write_request7_to_bank29   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank29    =  dma_read_addr7_to_bank29   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank29     =  read_request7_to_bank29    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank30
  wire dma_write_addr7_to_bank30      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr7_to_bank30       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank30   =  dma_write_addr7_to_bank30  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank30    =  write_request7_to_bank30   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank30    =  dma_read_addr7_to_bank30   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank30     =  read_request7_to_bank30    & memc__dma__read_ready7   ;                                         
  // DMA 7, bank31
  wire dma_write_addr7_to_bank31      =  (dma__memc__write_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr7_to_bank31       =  (dma__memc__read_address7[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank31   =  dma_write_addr7_to_bank31  & dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank31    =  write_request7_to_bank31   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank31    =  dma_read_addr7_to_bank31   & dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank31     =  read_request7_to_bank31    & memc__dma__read_ready7   ;                                         
  // DMA 8
  wire read_pause8     =  dma__memc__read_pause8   ;  
  // DMA 8, bank0
  wire dma_write_addr8_to_bank0      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr8_to_bank0       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank0   =  dma_write_addr8_to_bank0  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank0    =  write_request8_to_bank0   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank0    =  dma_read_addr8_to_bank0   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank0     =  read_request8_to_bank0    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank1
  wire dma_write_addr8_to_bank1      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr8_to_bank1       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank1   =  dma_write_addr8_to_bank1  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank1    =  write_request8_to_bank1   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank1    =  dma_read_addr8_to_bank1   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank1     =  read_request8_to_bank1    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank2
  wire dma_write_addr8_to_bank2      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr8_to_bank2       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank2   =  dma_write_addr8_to_bank2  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank2    =  write_request8_to_bank2   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank2    =  dma_read_addr8_to_bank2   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank2     =  read_request8_to_bank2    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank3
  wire dma_write_addr8_to_bank3      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr8_to_bank3       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank3   =  dma_write_addr8_to_bank3  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank3    =  write_request8_to_bank3   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank3    =  dma_read_addr8_to_bank3   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank3     =  read_request8_to_bank3    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank4
  wire dma_write_addr8_to_bank4      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr8_to_bank4       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank4   =  dma_write_addr8_to_bank4  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank4    =  write_request8_to_bank4   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank4    =  dma_read_addr8_to_bank4   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank4     =  read_request8_to_bank4    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank5
  wire dma_write_addr8_to_bank5      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr8_to_bank5       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank5   =  dma_write_addr8_to_bank5  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank5    =  write_request8_to_bank5   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank5    =  dma_read_addr8_to_bank5   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank5     =  read_request8_to_bank5    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank6
  wire dma_write_addr8_to_bank6      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr8_to_bank6       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank6   =  dma_write_addr8_to_bank6  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank6    =  write_request8_to_bank6   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank6    =  dma_read_addr8_to_bank6   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank6     =  read_request8_to_bank6    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank7
  wire dma_write_addr8_to_bank7      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr8_to_bank7       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank7   =  dma_write_addr8_to_bank7  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank7    =  write_request8_to_bank7   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank7    =  dma_read_addr8_to_bank7   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank7     =  read_request8_to_bank7    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank8
  wire dma_write_addr8_to_bank8      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr8_to_bank8       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank8   =  dma_write_addr8_to_bank8  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank8    =  write_request8_to_bank8   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank8    =  dma_read_addr8_to_bank8   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank8     =  read_request8_to_bank8    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank9
  wire dma_write_addr8_to_bank9      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr8_to_bank9       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank9   =  dma_write_addr8_to_bank9  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank9    =  write_request8_to_bank9   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank9    =  dma_read_addr8_to_bank9   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank9     =  read_request8_to_bank9    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank10
  wire dma_write_addr8_to_bank10      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr8_to_bank10       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank10   =  dma_write_addr8_to_bank10  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank10    =  write_request8_to_bank10   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank10    =  dma_read_addr8_to_bank10   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank10     =  read_request8_to_bank10    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank11
  wire dma_write_addr8_to_bank11      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr8_to_bank11       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank11   =  dma_write_addr8_to_bank11  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank11    =  write_request8_to_bank11   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank11    =  dma_read_addr8_to_bank11   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank11     =  read_request8_to_bank11    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank12
  wire dma_write_addr8_to_bank12      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr8_to_bank12       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank12   =  dma_write_addr8_to_bank12  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank12    =  write_request8_to_bank12   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank12    =  dma_read_addr8_to_bank12   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank12     =  read_request8_to_bank12    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank13
  wire dma_write_addr8_to_bank13      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr8_to_bank13       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank13   =  dma_write_addr8_to_bank13  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank13    =  write_request8_to_bank13   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank13    =  dma_read_addr8_to_bank13   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank13     =  read_request8_to_bank13    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank14
  wire dma_write_addr8_to_bank14      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr8_to_bank14       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank14   =  dma_write_addr8_to_bank14  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank14    =  write_request8_to_bank14   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank14    =  dma_read_addr8_to_bank14   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank14     =  read_request8_to_bank14    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank15
  wire dma_write_addr8_to_bank15      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr8_to_bank15       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank15   =  dma_write_addr8_to_bank15  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank15    =  write_request8_to_bank15   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank15    =  dma_read_addr8_to_bank15   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank15     =  read_request8_to_bank15    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank16
  wire dma_write_addr8_to_bank16      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr8_to_bank16       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank16   =  dma_write_addr8_to_bank16  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank16    =  write_request8_to_bank16   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank16    =  dma_read_addr8_to_bank16   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank16     =  read_request8_to_bank16    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank17
  wire dma_write_addr8_to_bank17      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr8_to_bank17       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank17   =  dma_write_addr8_to_bank17  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank17    =  write_request8_to_bank17   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank17    =  dma_read_addr8_to_bank17   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank17     =  read_request8_to_bank17    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank18
  wire dma_write_addr8_to_bank18      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr8_to_bank18       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank18   =  dma_write_addr8_to_bank18  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank18    =  write_request8_to_bank18   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank18    =  dma_read_addr8_to_bank18   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank18     =  read_request8_to_bank18    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank19
  wire dma_write_addr8_to_bank19      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr8_to_bank19       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank19   =  dma_write_addr8_to_bank19  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank19    =  write_request8_to_bank19   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank19    =  dma_read_addr8_to_bank19   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank19     =  read_request8_to_bank19    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank20
  wire dma_write_addr8_to_bank20      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr8_to_bank20       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank20   =  dma_write_addr8_to_bank20  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank20    =  write_request8_to_bank20   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank20    =  dma_read_addr8_to_bank20   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank20     =  read_request8_to_bank20    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank21
  wire dma_write_addr8_to_bank21      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr8_to_bank21       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank21   =  dma_write_addr8_to_bank21  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank21    =  write_request8_to_bank21   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank21    =  dma_read_addr8_to_bank21   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank21     =  read_request8_to_bank21    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank22
  wire dma_write_addr8_to_bank22      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr8_to_bank22       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank22   =  dma_write_addr8_to_bank22  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank22    =  write_request8_to_bank22   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank22    =  dma_read_addr8_to_bank22   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank22     =  read_request8_to_bank22    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank23
  wire dma_write_addr8_to_bank23      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr8_to_bank23       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank23   =  dma_write_addr8_to_bank23  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank23    =  write_request8_to_bank23   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank23    =  dma_read_addr8_to_bank23   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank23     =  read_request8_to_bank23    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank24
  wire dma_write_addr8_to_bank24      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr8_to_bank24       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank24   =  dma_write_addr8_to_bank24  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank24    =  write_request8_to_bank24   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank24    =  dma_read_addr8_to_bank24   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank24     =  read_request8_to_bank24    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank25
  wire dma_write_addr8_to_bank25      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr8_to_bank25       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank25   =  dma_write_addr8_to_bank25  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank25    =  write_request8_to_bank25   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank25    =  dma_read_addr8_to_bank25   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank25     =  read_request8_to_bank25    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank26
  wire dma_write_addr8_to_bank26      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr8_to_bank26       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank26   =  dma_write_addr8_to_bank26  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank26    =  write_request8_to_bank26   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank26    =  dma_read_addr8_to_bank26   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank26     =  read_request8_to_bank26    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank27
  wire dma_write_addr8_to_bank27      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr8_to_bank27       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank27   =  dma_write_addr8_to_bank27  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank27    =  write_request8_to_bank27   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank27    =  dma_read_addr8_to_bank27   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank27     =  read_request8_to_bank27    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank28
  wire dma_write_addr8_to_bank28      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr8_to_bank28       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank28   =  dma_write_addr8_to_bank28  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank28    =  write_request8_to_bank28   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank28    =  dma_read_addr8_to_bank28   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank28     =  read_request8_to_bank28    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank29
  wire dma_write_addr8_to_bank29      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr8_to_bank29       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank29   =  dma_write_addr8_to_bank29  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank29    =  write_request8_to_bank29   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank29    =  dma_read_addr8_to_bank29   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank29     =  read_request8_to_bank29    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank30
  wire dma_write_addr8_to_bank30      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr8_to_bank30       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank30   =  dma_write_addr8_to_bank30  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank30    =  write_request8_to_bank30   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank30    =  dma_read_addr8_to_bank30   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank30     =  read_request8_to_bank30    & memc__dma__read_ready8   ;                                         
  // DMA 8, bank31
  wire dma_write_addr8_to_bank31      =  (dma__memc__write_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr8_to_bank31       =  (dma__memc__read_address8[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank31   =  dma_write_addr8_to_bank31  & dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank31    =  write_request8_to_bank31   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank31    =  dma_read_addr8_to_bank31   & dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank31     =  read_request8_to_bank31    & memc__dma__read_ready8   ;                                         
  // DMA 9
  wire read_pause9     =  dma__memc__read_pause9   ;  
  // DMA 9, bank0
  wire dma_write_addr9_to_bank0      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr9_to_bank0       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank0   =  dma_write_addr9_to_bank0  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank0    =  write_request9_to_bank0   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank0    =  dma_read_addr9_to_bank0   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank0     =  read_request9_to_bank0    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank1
  wire dma_write_addr9_to_bank1      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr9_to_bank1       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank1   =  dma_write_addr9_to_bank1  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank1    =  write_request9_to_bank1   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank1    =  dma_read_addr9_to_bank1   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank1     =  read_request9_to_bank1    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank2
  wire dma_write_addr9_to_bank2      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr9_to_bank2       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank2   =  dma_write_addr9_to_bank2  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank2    =  write_request9_to_bank2   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank2    =  dma_read_addr9_to_bank2   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank2     =  read_request9_to_bank2    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank3
  wire dma_write_addr9_to_bank3      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr9_to_bank3       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank3   =  dma_write_addr9_to_bank3  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank3    =  write_request9_to_bank3   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank3    =  dma_read_addr9_to_bank3   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank3     =  read_request9_to_bank3    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank4
  wire dma_write_addr9_to_bank4      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr9_to_bank4       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank4   =  dma_write_addr9_to_bank4  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank4    =  write_request9_to_bank4   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank4    =  dma_read_addr9_to_bank4   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank4     =  read_request9_to_bank4    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank5
  wire dma_write_addr9_to_bank5      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr9_to_bank5       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank5   =  dma_write_addr9_to_bank5  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank5    =  write_request9_to_bank5   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank5    =  dma_read_addr9_to_bank5   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank5     =  read_request9_to_bank5    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank6
  wire dma_write_addr9_to_bank6      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr9_to_bank6       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank6   =  dma_write_addr9_to_bank6  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank6    =  write_request9_to_bank6   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank6    =  dma_read_addr9_to_bank6   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank6     =  read_request9_to_bank6    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank7
  wire dma_write_addr9_to_bank7      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr9_to_bank7       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank7   =  dma_write_addr9_to_bank7  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank7    =  write_request9_to_bank7   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank7    =  dma_read_addr9_to_bank7   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank7     =  read_request9_to_bank7    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank8
  wire dma_write_addr9_to_bank8      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr9_to_bank8       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank8   =  dma_write_addr9_to_bank8  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank8    =  write_request9_to_bank8   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank8    =  dma_read_addr9_to_bank8   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank8     =  read_request9_to_bank8    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank9
  wire dma_write_addr9_to_bank9      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr9_to_bank9       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank9   =  dma_write_addr9_to_bank9  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank9    =  write_request9_to_bank9   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank9    =  dma_read_addr9_to_bank9   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank9     =  read_request9_to_bank9    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank10
  wire dma_write_addr9_to_bank10      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr9_to_bank10       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank10   =  dma_write_addr9_to_bank10  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank10    =  write_request9_to_bank10   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank10    =  dma_read_addr9_to_bank10   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank10     =  read_request9_to_bank10    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank11
  wire dma_write_addr9_to_bank11      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr9_to_bank11       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank11   =  dma_write_addr9_to_bank11  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank11    =  write_request9_to_bank11   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank11    =  dma_read_addr9_to_bank11   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank11     =  read_request9_to_bank11    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank12
  wire dma_write_addr9_to_bank12      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr9_to_bank12       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank12   =  dma_write_addr9_to_bank12  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank12    =  write_request9_to_bank12   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank12    =  dma_read_addr9_to_bank12   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank12     =  read_request9_to_bank12    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank13
  wire dma_write_addr9_to_bank13      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr9_to_bank13       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank13   =  dma_write_addr9_to_bank13  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank13    =  write_request9_to_bank13   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank13    =  dma_read_addr9_to_bank13   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank13     =  read_request9_to_bank13    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank14
  wire dma_write_addr9_to_bank14      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr9_to_bank14       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank14   =  dma_write_addr9_to_bank14  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank14    =  write_request9_to_bank14   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank14    =  dma_read_addr9_to_bank14   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank14     =  read_request9_to_bank14    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank15
  wire dma_write_addr9_to_bank15      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr9_to_bank15       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank15   =  dma_write_addr9_to_bank15  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank15    =  write_request9_to_bank15   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank15    =  dma_read_addr9_to_bank15   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank15     =  read_request9_to_bank15    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank16
  wire dma_write_addr9_to_bank16      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr9_to_bank16       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank16   =  dma_write_addr9_to_bank16  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank16    =  write_request9_to_bank16   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank16    =  dma_read_addr9_to_bank16   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank16     =  read_request9_to_bank16    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank17
  wire dma_write_addr9_to_bank17      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr9_to_bank17       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank17   =  dma_write_addr9_to_bank17  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank17    =  write_request9_to_bank17   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank17    =  dma_read_addr9_to_bank17   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank17     =  read_request9_to_bank17    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank18
  wire dma_write_addr9_to_bank18      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr9_to_bank18       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank18   =  dma_write_addr9_to_bank18  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank18    =  write_request9_to_bank18   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank18    =  dma_read_addr9_to_bank18   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank18     =  read_request9_to_bank18    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank19
  wire dma_write_addr9_to_bank19      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr9_to_bank19       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank19   =  dma_write_addr9_to_bank19  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank19    =  write_request9_to_bank19   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank19    =  dma_read_addr9_to_bank19   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank19     =  read_request9_to_bank19    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank20
  wire dma_write_addr9_to_bank20      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr9_to_bank20       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank20   =  dma_write_addr9_to_bank20  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank20    =  write_request9_to_bank20   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank20    =  dma_read_addr9_to_bank20   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank20     =  read_request9_to_bank20    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank21
  wire dma_write_addr9_to_bank21      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr9_to_bank21       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank21   =  dma_write_addr9_to_bank21  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank21    =  write_request9_to_bank21   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank21    =  dma_read_addr9_to_bank21   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank21     =  read_request9_to_bank21    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank22
  wire dma_write_addr9_to_bank22      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr9_to_bank22       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank22   =  dma_write_addr9_to_bank22  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank22    =  write_request9_to_bank22   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank22    =  dma_read_addr9_to_bank22   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank22     =  read_request9_to_bank22    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank23
  wire dma_write_addr9_to_bank23      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr9_to_bank23       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank23   =  dma_write_addr9_to_bank23  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank23    =  write_request9_to_bank23   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank23    =  dma_read_addr9_to_bank23   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank23     =  read_request9_to_bank23    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank24
  wire dma_write_addr9_to_bank24      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr9_to_bank24       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank24   =  dma_write_addr9_to_bank24  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank24    =  write_request9_to_bank24   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank24    =  dma_read_addr9_to_bank24   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank24     =  read_request9_to_bank24    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank25
  wire dma_write_addr9_to_bank25      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr9_to_bank25       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank25   =  dma_write_addr9_to_bank25  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank25    =  write_request9_to_bank25   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank25    =  dma_read_addr9_to_bank25   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank25     =  read_request9_to_bank25    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank26
  wire dma_write_addr9_to_bank26      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr9_to_bank26       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank26   =  dma_write_addr9_to_bank26  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank26    =  write_request9_to_bank26   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank26    =  dma_read_addr9_to_bank26   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank26     =  read_request9_to_bank26    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank27
  wire dma_write_addr9_to_bank27      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr9_to_bank27       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank27   =  dma_write_addr9_to_bank27  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank27    =  write_request9_to_bank27   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank27    =  dma_read_addr9_to_bank27   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank27     =  read_request9_to_bank27    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank28
  wire dma_write_addr9_to_bank28      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr9_to_bank28       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank28   =  dma_write_addr9_to_bank28  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank28    =  write_request9_to_bank28   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank28    =  dma_read_addr9_to_bank28   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank28     =  read_request9_to_bank28    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank29
  wire dma_write_addr9_to_bank29      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr9_to_bank29       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank29   =  dma_write_addr9_to_bank29  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank29    =  write_request9_to_bank29   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank29    =  dma_read_addr9_to_bank29   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank29     =  read_request9_to_bank29    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank30
  wire dma_write_addr9_to_bank30      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr9_to_bank30       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank30   =  dma_write_addr9_to_bank30  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank30    =  write_request9_to_bank30   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank30    =  dma_read_addr9_to_bank30   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank30     =  read_request9_to_bank30    & memc__dma__read_ready9   ;                                         
  // DMA 9, bank31
  wire dma_write_addr9_to_bank31      =  (dma__memc__write_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr9_to_bank31       =  (dma__memc__read_address9[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank31   =  dma_write_addr9_to_bank31  & dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank31    =  write_request9_to_bank31   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank31    =  dma_read_addr9_to_bank31   & dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank31     =  read_request9_to_bank31    & memc__dma__read_ready9   ;                                         
  // DMA 10
  wire read_pause10     =  dma__memc__read_pause10   ;  
  // DMA 10, bank0
  wire dma_write_addr10_to_bank0      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr10_to_bank0       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank0   =  dma_write_addr10_to_bank0  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank0    =  write_request10_to_bank0   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank0    =  dma_read_addr10_to_bank0   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank0     =  read_request10_to_bank0    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank1
  wire dma_write_addr10_to_bank1      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr10_to_bank1       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank1   =  dma_write_addr10_to_bank1  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank1    =  write_request10_to_bank1   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank1    =  dma_read_addr10_to_bank1   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank1     =  read_request10_to_bank1    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank2
  wire dma_write_addr10_to_bank2      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr10_to_bank2       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank2   =  dma_write_addr10_to_bank2  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank2    =  write_request10_to_bank2   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank2    =  dma_read_addr10_to_bank2   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank2     =  read_request10_to_bank2    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank3
  wire dma_write_addr10_to_bank3      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr10_to_bank3       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank3   =  dma_write_addr10_to_bank3  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank3    =  write_request10_to_bank3   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank3    =  dma_read_addr10_to_bank3   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank3     =  read_request10_to_bank3    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank4
  wire dma_write_addr10_to_bank4      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr10_to_bank4       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank4   =  dma_write_addr10_to_bank4  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank4    =  write_request10_to_bank4   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank4    =  dma_read_addr10_to_bank4   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank4     =  read_request10_to_bank4    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank5
  wire dma_write_addr10_to_bank5      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr10_to_bank5       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank5   =  dma_write_addr10_to_bank5  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank5    =  write_request10_to_bank5   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank5    =  dma_read_addr10_to_bank5   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank5     =  read_request10_to_bank5    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank6
  wire dma_write_addr10_to_bank6      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr10_to_bank6       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank6   =  dma_write_addr10_to_bank6  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank6    =  write_request10_to_bank6   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank6    =  dma_read_addr10_to_bank6   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank6     =  read_request10_to_bank6    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank7
  wire dma_write_addr10_to_bank7      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr10_to_bank7       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank7   =  dma_write_addr10_to_bank7  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank7    =  write_request10_to_bank7   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank7    =  dma_read_addr10_to_bank7   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank7     =  read_request10_to_bank7    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank8
  wire dma_write_addr10_to_bank8      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr10_to_bank8       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank8   =  dma_write_addr10_to_bank8  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank8    =  write_request10_to_bank8   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank8    =  dma_read_addr10_to_bank8   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank8     =  read_request10_to_bank8    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank9
  wire dma_write_addr10_to_bank9      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr10_to_bank9       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank9   =  dma_write_addr10_to_bank9  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank9    =  write_request10_to_bank9   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank9    =  dma_read_addr10_to_bank9   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank9     =  read_request10_to_bank9    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank10
  wire dma_write_addr10_to_bank10      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr10_to_bank10       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank10   =  dma_write_addr10_to_bank10  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank10    =  write_request10_to_bank10   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank10    =  dma_read_addr10_to_bank10   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank10     =  read_request10_to_bank10    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank11
  wire dma_write_addr10_to_bank11      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr10_to_bank11       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank11   =  dma_write_addr10_to_bank11  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank11    =  write_request10_to_bank11   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank11    =  dma_read_addr10_to_bank11   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank11     =  read_request10_to_bank11    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank12
  wire dma_write_addr10_to_bank12      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr10_to_bank12       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank12   =  dma_write_addr10_to_bank12  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank12    =  write_request10_to_bank12   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank12    =  dma_read_addr10_to_bank12   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank12     =  read_request10_to_bank12    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank13
  wire dma_write_addr10_to_bank13      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr10_to_bank13       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank13   =  dma_write_addr10_to_bank13  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank13    =  write_request10_to_bank13   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank13    =  dma_read_addr10_to_bank13   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank13     =  read_request10_to_bank13    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank14
  wire dma_write_addr10_to_bank14      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr10_to_bank14       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank14   =  dma_write_addr10_to_bank14  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank14    =  write_request10_to_bank14   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank14    =  dma_read_addr10_to_bank14   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank14     =  read_request10_to_bank14    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank15
  wire dma_write_addr10_to_bank15      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr10_to_bank15       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank15   =  dma_write_addr10_to_bank15  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank15    =  write_request10_to_bank15   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank15    =  dma_read_addr10_to_bank15   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank15     =  read_request10_to_bank15    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank16
  wire dma_write_addr10_to_bank16      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr10_to_bank16       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank16   =  dma_write_addr10_to_bank16  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank16    =  write_request10_to_bank16   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank16    =  dma_read_addr10_to_bank16   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank16     =  read_request10_to_bank16    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank17
  wire dma_write_addr10_to_bank17      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr10_to_bank17       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank17   =  dma_write_addr10_to_bank17  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank17    =  write_request10_to_bank17   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank17    =  dma_read_addr10_to_bank17   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank17     =  read_request10_to_bank17    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank18
  wire dma_write_addr10_to_bank18      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr10_to_bank18       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank18   =  dma_write_addr10_to_bank18  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank18    =  write_request10_to_bank18   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank18    =  dma_read_addr10_to_bank18   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank18     =  read_request10_to_bank18    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank19
  wire dma_write_addr10_to_bank19      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr10_to_bank19       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank19   =  dma_write_addr10_to_bank19  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank19    =  write_request10_to_bank19   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank19    =  dma_read_addr10_to_bank19   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank19     =  read_request10_to_bank19    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank20
  wire dma_write_addr10_to_bank20      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr10_to_bank20       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank20   =  dma_write_addr10_to_bank20  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank20    =  write_request10_to_bank20   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank20    =  dma_read_addr10_to_bank20   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank20     =  read_request10_to_bank20    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank21
  wire dma_write_addr10_to_bank21      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr10_to_bank21       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank21   =  dma_write_addr10_to_bank21  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank21    =  write_request10_to_bank21   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank21    =  dma_read_addr10_to_bank21   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank21     =  read_request10_to_bank21    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank22
  wire dma_write_addr10_to_bank22      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr10_to_bank22       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank22   =  dma_write_addr10_to_bank22  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank22    =  write_request10_to_bank22   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank22    =  dma_read_addr10_to_bank22   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank22     =  read_request10_to_bank22    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank23
  wire dma_write_addr10_to_bank23      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr10_to_bank23       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank23   =  dma_write_addr10_to_bank23  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank23    =  write_request10_to_bank23   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank23    =  dma_read_addr10_to_bank23   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank23     =  read_request10_to_bank23    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank24
  wire dma_write_addr10_to_bank24      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr10_to_bank24       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank24   =  dma_write_addr10_to_bank24  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank24    =  write_request10_to_bank24   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank24    =  dma_read_addr10_to_bank24   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank24     =  read_request10_to_bank24    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank25
  wire dma_write_addr10_to_bank25      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr10_to_bank25       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank25   =  dma_write_addr10_to_bank25  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank25    =  write_request10_to_bank25   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank25    =  dma_read_addr10_to_bank25   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank25     =  read_request10_to_bank25    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank26
  wire dma_write_addr10_to_bank26      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr10_to_bank26       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank26   =  dma_write_addr10_to_bank26  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank26    =  write_request10_to_bank26   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank26    =  dma_read_addr10_to_bank26   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank26     =  read_request10_to_bank26    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank27
  wire dma_write_addr10_to_bank27      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr10_to_bank27       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank27   =  dma_write_addr10_to_bank27  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank27    =  write_request10_to_bank27   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank27    =  dma_read_addr10_to_bank27   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank27     =  read_request10_to_bank27    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank28
  wire dma_write_addr10_to_bank28      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr10_to_bank28       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank28   =  dma_write_addr10_to_bank28  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank28    =  write_request10_to_bank28   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank28    =  dma_read_addr10_to_bank28   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank28     =  read_request10_to_bank28    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank29
  wire dma_write_addr10_to_bank29      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr10_to_bank29       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank29   =  dma_write_addr10_to_bank29  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank29    =  write_request10_to_bank29   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank29    =  dma_read_addr10_to_bank29   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank29     =  read_request10_to_bank29    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank30
  wire dma_write_addr10_to_bank30      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr10_to_bank30       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank30   =  dma_write_addr10_to_bank30  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank30    =  write_request10_to_bank30   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank30    =  dma_read_addr10_to_bank30   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank30     =  read_request10_to_bank30    & memc__dma__read_ready10   ;                                         
  // DMA 10, bank31
  wire dma_write_addr10_to_bank31      =  (dma__memc__write_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr10_to_bank31       =  (dma__memc__read_address10[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank31   =  dma_write_addr10_to_bank31  & dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank31    =  write_request10_to_bank31   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank31    =  dma_read_addr10_to_bank31   & dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank31     =  read_request10_to_bank31    & memc__dma__read_ready10   ;                                         
  // DMA 11
  wire read_pause11     =  dma__memc__read_pause11   ;  
  // DMA 11, bank0
  wire dma_write_addr11_to_bank0      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr11_to_bank0       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank0   =  dma_write_addr11_to_bank0  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank0    =  write_request11_to_bank0   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank0    =  dma_read_addr11_to_bank0   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank0     =  read_request11_to_bank0    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank1
  wire dma_write_addr11_to_bank1      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr11_to_bank1       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank1   =  dma_write_addr11_to_bank1  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank1    =  write_request11_to_bank1   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank1    =  dma_read_addr11_to_bank1   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank1     =  read_request11_to_bank1    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank2
  wire dma_write_addr11_to_bank2      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr11_to_bank2       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank2   =  dma_write_addr11_to_bank2  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank2    =  write_request11_to_bank2   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank2    =  dma_read_addr11_to_bank2   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank2     =  read_request11_to_bank2    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank3
  wire dma_write_addr11_to_bank3      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr11_to_bank3       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank3   =  dma_write_addr11_to_bank3  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank3    =  write_request11_to_bank3   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank3    =  dma_read_addr11_to_bank3   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank3     =  read_request11_to_bank3    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank4
  wire dma_write_addr11_to_bank4      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr11_to_bank4       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank4   =  dma_write_addr11_to_bank4  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank4    =  write_request11_to_bank4   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank4    =  dma_read_addr11_to_bank4   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank4     =  read_request11_to_bank4    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank5
  wire dma_write_addr11_to_bank5      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr11_to_bank5       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank5   =  dma_write_addr11_to_bank5  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank5    =  write_request11_to_bank5   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank5    =  dma_read_addr11_to_bank5   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank5     =  read_request11_to_bank5    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank6
  wire dma_write_addr11_to_bank6      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr11_to_bank6       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank6   =  dma_write_addr11_to_bank6  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank6    =  write_request11_to_bank6   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank6    =  dma_read_addr11_to_bank6   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank6     =  read_request11_to_bank6    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank7
  wire dma_write_addr11_to_bank7      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr11_to_bank7       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank7   =  dma_write_addr11_to_bank7  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank7    =  write_request11_to_bank7   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank7    =  dma_read_addr11_to_bank7   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank7     =  read_request11_to_bank7    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank8
  wire dma_write_addr11_to_bank8      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr11_to_bank8       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank8   =  dma_write_addr11_to_bank8  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank8    =  write_request11_to_bank8   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank8    =  dma_read_addr11_to_bank8   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank8     =  read_request11_to_bank8    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank9
  wire dma_write_addr11_to_bank9      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr11_to_bank9       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank9   =  dma_write_addr11_to_bank9  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank9    =  write_request11_to_bank9   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank9    =  dma_read_addr11_to_bank9   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank9     =  read_request11_to_bank9    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank10
  wire dma_write_addr11_to_bank10      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr11_to_bank10       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank10   =  dma_write_addr11_to_bank10  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank10    =  write_request11_to_bank10   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank10    =  dma_read_addr11_to_bank10   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank10     =  read_request11_to_bank10    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank11
  wire dma_write_addr11_to_bank11      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr11_to_bank11       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank11   =  dma_write_addr11_to_bank11  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank11    =  write_request11_to_bank11   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank11    =  dma_read_addr11_to_bank11   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank11     =  read_request11_to_bank11    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank12
  wire dma_write_addr11_to_bank12      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr11_to_bank12       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank12   =  dma_write_addr11_to_bank12  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank12    =  write_request11_to_bank12   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank12    =  dma_read_addr11_to_bank12   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank12     =  read_request11_to_bank12    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank13
  wire dma_write_addr11_to_bank13      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr11_to_bank13       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank13   =  dma_write_addr11_to_bank13  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank13    =  write_request11_to_bank13   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank13    =  dma_read_addr11_to_bank13   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank13     =  read_request11_to_bank13    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank14
  wire dma_write_addr11_to_bank14      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr11_to_bank14       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank14   =  dma_write_addr11_to_bank14  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank14    =  write_request11_to_bank14   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank14    =  dma_read_addr11_to_bank14   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank14     =  read_request11_to_bank14    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank15
  wire dma_write_addr11_to_bank15      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr11_to_bank15       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank15   =  dma_write_addr11_to_bank15  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank15    =  write_request11_to_bank15   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank15    =  dma_read_addr11_to_bank15   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank15     =  read_request11_to_bank15    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank16
  wire dma_write_addr11_to_bank16      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr11_to_bank16       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank16   =  dma_write_addr11_to_bank16  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank16    =  write_request11_to_bank16   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank16    =  dma_read_addr11_to_bank16   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank16     =  read_request11_to_bank16    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank17
  wire dma_write_addr11_to_bank17      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr11_to_bank17       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank17   =  dma_write_addr11_to_bank17  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank17    =  write_request11_to_bank17   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank17    =  dma_read_addr11_to_bank17   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank17     =  read_request11_to_bank17    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank18
  wire dma_write_addr11_to_bank18      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr11_to_bank18       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank18   =  dma_write_addr11_to_bank18  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank18    =  write_request11_to_bank18   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank18    =  dma_read_addr11_to_bank18   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank18     =  read_request11_to_bank18    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank19
  wire dma_write_addr11_to_bank19      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr11_to_bank19       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank19   =  dma_write_addr11_to_bank19  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank19    =  write_request11_to_bank19   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank19    =  dma_read_addr11_to_bank19   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank19     =  read_request11_to_bank19    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank20
  wire dma_write_addr11_to_bank20      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr11_to_bank20       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank20   =  dma_write_addr11_to_bank20  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank20    =  write_request11_to_bank20   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank20    =  dma_read_addr11_to_bank20   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank20     =  read_request11_to_bank20    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank21
  wire dma_write_addr11_to_bank21      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr11_to_bank21       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank21   =  dma_write_addr11_to_bank21  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank21    =  write_request11_to_bank21   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank21    =  dma_read_addr11_to_bank21   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank21     =  read_request11_to_bank21    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank22
  wire dma_write_addr11_to_bank22      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr11_to_bank22       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank22   =  dma_write_addr11_to_bank22  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank22    =  write_request11_to_bank22   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank22    =  dma_read_addr11_to_bank22   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank22     =  read_request11_to_bank22    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank23
  wire dma_write_addr11_to_bank23      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr11_to_bank23       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank23   =  dma_write_addr11_to_bank23  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank23    =  write_request11_to_bank23   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank23    =  dma_read_addr11_to_bank23   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank23     =  read_request11_to_bank23    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank24
  wire dma_write_addr11_to_bank24      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr11_to_bank24       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank24   =  dma_write_addr11_to_bank24  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank24    =  write_request11_to_bank24   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank24    =  dma_read_addr11_to_bank24   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank24     =  read_request11_to_bank24    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank25
  wire dma_write_addr11_to_bank25      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr11_to_bank25       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank25   =  dma_write_addr11_to_bank25  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank25    =  write_request11_to_bank25   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank25    =  dma_read_addr11_to_bank25   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank25     =  read_request11_to_bank25    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank26
  wire dma_write_addr11_to_bank26      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr11_to_bank26       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank26   =  dma_write_addr11_to_bank26  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank26    =  write_request11_to_bank26   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank26    =  dma_read_addr11_to_bank26   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank26     =  read_request11_to_bank26    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank27
  wire dma_write_addr11_to_bank27      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr11_to_bank27       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank27   =  dma_write_addr11_to_bank27  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank27    =  write_request11_to_bank27   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank27    =  dma_read_addr11_to_bank27   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank27     =  read_request11_to_bank27    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank28
  wire dma_write_addr11_to_bank28      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr11_to_bank28       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank28   =  dma_write_addr11_to_bank28  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank28    =  write_request11_to_bank28   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank28    =  dma_read_addr11_to_bank28   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank28     =  read_request11_to_bank28    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank29
  wire dma_write_addr11_to_bank29      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr11_to_bank29       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank29   =  dma_write_addr11_to_bank29  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank29    =  write_request11_to_bank29   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank29    =  dma_read_addr11_to_bank29   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank29     =  read_request11_to_bank29    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank30
  wire dma_write_addr11_to_bank30      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr11_to_bank30       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank30   =  dma_write_addr11_to_bank30  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank30    =  write_request11_to_bank30   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank30    =  dma_read_addr11_to_bank30   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank30     =  read_request11_to_bank30    & memc__dma__read_ready11   ;                                         
  // DMA 11, bank31
  wire dma_write_addr11_to_bank31      =  (dma__memc__write_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr11_to_bank31       =  (dma__memc__read_address11[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank31   =  dma_write_addr11_to_bank31  & dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank31    =  write_request11_to_bank31   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank31    =  dma_read_addr11_to_bank31   & dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank31     =  read_request11_to_bank31    & memc__dma__read_ready11   ;                                         
  // DMA 12
  wire read_pause12     =  dma__memc__read_pause12   ;  
  // DMA 12, bank0
  wire dma_write_addr12_to_bank0      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr12_to_bank0       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank0   =  dma_write_addr12_to_bank0  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank0    =  write_request12_to_bank0   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank0    =  dma_read_addr12_to_bank0   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank0     =  read_request12_to_bank0    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank1
  wire dma_write_addr12_to_bank1      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr12_to_bank1       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank1   =  dma_write_addr12_to_bank1  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank1    =  write_request12_to_bank1   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank1    =  dma_read_addr12_to_bank1   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank1     =  read_request12_to_bank1    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank2
  wire dma_write_addr12_to_bank2      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr12_to_bank2       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank2   =  dma_write_addr12_to_bank2  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank2    =  write_request12_to_bank2   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank2    =  dma_read_addr12_to_bank2   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank2     =  read_request12_to_bank2    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank3
  wire dma_write_addr12_to_bank3      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr12_to_bank3       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank3   =  dma_write_addr12_to_bank3  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank3    =  write_request12_to_bank3   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank3    =  dma_read_addr12_to_bank3   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank3     =  read_request12_to_bank3    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank4
  wire dma_write_addr12_to_bank4      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr12_to_bank4       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank4   =  dma_write_addr12_to_bank4  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank4    =  write_request12_to_bank4   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank4    =  dma_read_addr12_to_bank4   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank4     =  read_request12_to_bank4    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank5
  wire dma_write_addr12_to_bank5      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr12_to_bank5       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank5   =  dma_write_addr12_to_bank5  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank5    =  write_request12_to_bank5   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank5    =  dma_read_addr12_to_bank5   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank5     =  read_request12_to_bank5    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank6
  wire dma_write_addr12_to_bank6      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr12_to_bank6       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank6   =  dma_write_addr12_to_bank6  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank6    =  write_request12_to_bank6   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank6    =  dma_read_addr12_to_bank6   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank6     =  read_request12_to_bank6    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank7
  wire dma_write_addr12_to_bank7      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr12_to_bank7       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank7   =  dma_write_addr12_to_bank7  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank7    =  write_request12_to_bank7   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank7    =  dma_read_addr12_to_bank7   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank7     =  read_request12_to_bank7    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank8
  wire dma_write_addr12_to_bank8      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr12_to_bank8       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank8   =  dma_write_addr12_to_bank8  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank8    =  write_request12_to_bank8   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank8    =  dma_read_addr12_to_bank8   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank8     =  read_request12_to_bank8    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank9
  wire dma_write_addr12_to_bank9      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr12_to_bank9       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank9   =  dma_write_addr12_to_bank9  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank9    =  write_request12_to_bank9   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank9    =  dma_read_addr12_to_bank9   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank9     =  read_request12_to_bank9    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank10
  wire dma_write_addr12_to_bank10      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr12_to_bank10       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank10   =  dma_write_addr12_to_bank10  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank10    =  write_request12_to_bank10   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank10    =  dma_read_addr12_to_bank10   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank10     =  read_request12_to_bank10    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank11
  wire dma_write_addr12_to_bank11      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr12_to_bank11       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank11   =  dma_write_addr12_to_bank11  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank11    =  write_request12_to_bank11   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank11    =  dma_read_addr12_to_bank11   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank11     =  read_request12_to_bank11    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank12
  wire dma_write_addr12_to_bank12      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr12_to_bank12       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank12   =  dma_write_addr12_to_bank12  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank12    =  write_request12_to_bank12   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank12    =  dma_read_addr12_to_bank12   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank12     =  read_request12_to_bank12    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank13
  wire dma_write_addr12_to_bank13      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr12_to_bank13       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank13   =  dma_write_addr12_to_bank13  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank13    =  write_request12_to_bank13   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank13    =  dma_read_addr12_to_bank13   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank13     =  read_request12_to_bank13    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank14
  wire dma_write_addr12_to_bank14      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr12_to_bank14       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank14   =  dma_write_addr12_to_bank14  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank14    =  write_request12_to_bank14   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank14    =  dma_read_addr12_to_bank14   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank14     =  read_request12_to_bank14    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank15
  wire dma_write_addr12_to_bank15      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr12_to_bank15       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank15   =  dma_write_addr12_to_bank15  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank15    =  write_request12_to_bank15   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank15    =  dma_read_addr12_to_bank15   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank15     =  read_request12_to_bank15    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank16
  wire dma_write_addr12_to_bank16      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr12_to_bank16       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank16   =  dma_write_addr12_to_bank16  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank16    =  write_request12_to_bank16   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank16    =  dma_read_addr12_to_bank16   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank16     =  read_request12_to_bank16    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank17
  wire dma_write_addr12_to_bank17      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr12_to_bank17       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank17   =  dma_write_addr12_to_bank17  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank17    =  write_request12_to_bank17   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank17    =  dma_read_addr12_to_bank17   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank17     =  read_request12_to_bank17    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank18
  wire dma_write_addr12_to_bank18      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr12_to_bank18       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank18   =  dma_write_addr12_to_bank18  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank18    =  write_request12_to_bank18   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank18    =  dma_read_addr12_to_bank18   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank18     =  read_request12_to_bank18    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank19
  wire dma_write_addr12_to_bank19      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr12_to_bank19       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank19   =  dma_write_addr12_to_bank19  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank19    =  write_request12_to_bank19   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank19    =  dma_read_addr12_to_bank19   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank19     =  read_request12_to_bank19    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank20
  wire dma_write_addr12_to_bank20      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr12_to_bank20       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank20   =  dma_write_addr12_to_bank20  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank20    =  write_request12_to_bank20   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank20    =  dma_read_addr12_to_bank20   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank20     =  read_request12_to_bank20    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank21
  wire dma_write_addr12_to_bank21      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr12_to_bank21       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank21   =  dma_write_addr12_to_bank21  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank21    =  write_request12_to_bank21   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank21    =  dma_read_addr12_to_bank21   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank21     =  read_request12_to_bank21    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank22
  wire dma_write_addr12_to_bank22      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr12_to_bank22       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank22   =  dma_write_addr12_to_bank22  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank22    =  write_request12_to_bank22   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank22    =  dma_read_addr12_to_bank22   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank22     =  read_request12_to_bank22    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank23
  wire dma_write_addr12_to_bank23      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr12_to_bank23       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank23   =  dma_write_addr12_to_bank23  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank23    =  write_request12_to_bank23   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank23    =  dma_read_addr12_to_bank23   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank23     =  read_request12_to_bank23    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank24
  wire dma_write_addr12_to_bank24      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr12_to_bank24       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank24   =  dma_write_addr12_to_bank24  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank24    =  write_request12_to_bank24   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank24    =  dma_read_addr12_to_bank24   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank24     =  read_request12_to_bank24    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank25
  wire dma_write_addr12_to_bank25      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr12_to_bank25       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank25   =  dma_write_addr12_to_bank25  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank25    =  write_request12_to_bank25   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank25    =  dma_read_addr12_to_bank25   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank25     =  read_request12_to_bank25    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank26
  wire dma_write_addr12_to_bank26      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr12_to_bank26       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank26   =  dma_write_addr12_to_bank26  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank26    =  write_request12_to_bank26   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank26    =  dma_read_addr12_to_bank26   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank26     =  read_request12_to_bank26    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank27
  wire dma_write_addr12_to_bank27      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr12_to_bank27       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank27   =  dma_write_addr12_to_bank27  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank27    =  write_request12_to_bank27   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank27    =  dma_read_addr12_to_bank27   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank27     =  read_request12_to_bank27    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank28
  wire dma_write_addr12_to_bank28      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr12_to_bank28       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank28   =  dma_write_addr12_to_bank28  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank28    =  write_request12_to_bank28   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank28    =  dma_read_addr12_to_bank28   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank28     =  read_request12_to_bank28    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank29
  wire dma_write_addr12_to_bank29      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr12_to_bank29       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank29   =  dma_write_addr12_to_bank29  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank29    =  write_request12_to_bank29   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank29    =  dma_read_addr12_to_bank29   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank29     =  read_request12_to_bank29    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank30
  wire dma_write_addr12_to_bank30      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr12_to_bank30       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank30   =  dma_write_addr12_to_bank30  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank30    =  write_request12_to_bank30   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank30    =  dma_read_addr12_to_bank30   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank30     =  read_request12_to_bank30    & memc__dma__read_ready12   ;                                         
  // DMA 12, bank31
  wire dma_write_addr12_to_bank31      =  (dma__memc__write_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr12_to_bank31       =  (dma__memc__read_address12[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank31   =  dma_write_addr12_to_bank31  & dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank31    =  write_request12_to_bank31   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank31    =  dma_read_addr12_to_bank31   & dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank31     =  read_request12_to_bank31    & memc__dma__read_ready12   ;                                         
  // DMA 13
  wire read_pause13     =  dma__memc__read_pause13   ;  
  // DMA 13, bank0
  wire dma_write_addr13_to_bank0      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr13_to_bank0       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank0   =  dma_write_addr13_to_bank0  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank0    =  write_request13_to_bank0   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank0    =  dma_read_addr13_to_bank0   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank0     =  read_request13_to_bank0    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank1
  wire dma_write_addr13_to_bank1      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr13_to_bank1       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank1   =  dma_write_addr13_to_bank1  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank1    =  write_request13_to_bank1   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank1    =  dma_read_addr13_to_bank1   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank1     =  read_request13_to_bank1    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank2
  wire dma_write_addr13_to_bank2      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr13_to_bank2       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank2   =  dma_write_addr13_to_bank2  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank2    =  write_request13_to_bank2   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank2    =  dma_read_addr13_to_bank2   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank2     =  read_request13_to_bank2    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank3
  wire dma_write_addr13_to_bank3      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr13_to_bank3       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank3   =  dma_write_addr13_to_bank3  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank3    =  write_request13_to_bank3   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank3    =  dma_read_addr13_to_bank3   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank3     =  read_request13_to_bank3    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank4
  wire dma_write_addr13_to_bank4      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr13_to_bank4       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank4   =  dma_write_addr13_to_bank4  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank4    =  write_request13_to_bank4   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank4    =  dma_read_addr13_to_bank4   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank4     =  read_request13_to_bank4    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank5
  wire dma_write_addr13_to_bank5      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr13_to_bank5       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank5   =  dma_write_addr13_to_bank5  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank5    =  write_request13_to_bank5   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank5    =  dma_read_addr13_to_bank5   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank5     =  read_request13_to_bank5    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank6
  wire dma_write_addr13_to_bank6      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr13_to_bank6       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank6   =  dma_write_addr13_to_bank6  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank6    =  write_request13_to_bank6   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank6    =  dma_read_addr13_to_bank6   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank6     =  read_request13_to_bank6    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank7
  wire dma_write_addr13_to_bank7      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr13_to_bank7       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank7   =  dma_write_addr13_to_bank7  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank7    =  write_request13_to_bank7   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank7    =  dma_read_addr13_to_bank7   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank7     =  read_request13_to_bank7    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank8
  wire dma_write_addr13_to_bank8      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr13_to_bank8       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank8   =  dma_write_addr13_to_bank8  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank8    =  write_request13_to_bank8   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank8    =  dma_read_addr13_to_bank8   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank8     =  read_request13_to_bank8    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank9
  wire dma_write_addr13_to_bank9      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr13_to_bank9       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank9   =  dma_write_addr13_to_bank9  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank9    =  write_request13_to_bank9   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank9    =  dma_read_addr13_to_bank9   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank9     =  read_request13_to_bank9    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank10
  wire dma_write_addr13_to_bank10      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr13_to_bank10       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank10   =  dma_write_addr13_to_bank10  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank10    =  write_request13_to_bank10   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank10    =  dma_read_addr13_to_bank10   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank10     =  read_request13_to_bank10    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank11
  wire dma_write_addr13_to_bank11      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr13_to_bank11       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank11   =  dma_write_addr13_to_bank11  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank11    =  write_request13_to_bank11   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank11    =  dma_read_addr13_to_bank11   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank11     =  read_request13_to_bank11    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank12
  wire dma_write_addr13_to_bank12      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr13_to_bank12       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank12   =  dma_write_addr13_to_bank12  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank12    =  write_request13_to_bank12   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank12    =  dma_read_addr13_to_bank12   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank12     =  read_request13_to_bank12    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank13
  wire dma_write_addr13_to_bank13      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr13_to_bank13       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank13   =  dma_write_addr13_to_bank13  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank13    =  write_request13_to_bank13   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank13    =  dma_read_addr13_to_bank13   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank13     =  read_request13_to_bank13    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank14
  wire dma_write_addr13_to_bank14      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr13_to_bank14       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank14   =  dma_write_addr13_to_bank14  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank14    =  write_request13_to_bank14   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank14    =  dma_read_addr13_to_bank14   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank14     =  read_request13_to_bank14    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank15
  wire dma_write_addr13_to_bank15      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr13_to_bank15       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank15   =  dma_write_addr13_to_bank15  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank15    =  write_request13_to_bank15   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank15    =  dma_read_addr13_to_bank15   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank15     =  read_request13_to_bank15    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank16
  wire dma_write_addr13_to_bank16      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr13_to_bank16       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank16   =  dma_write_addr13_to_bank16  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank16    =  write_request13_to_bank16   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank16    =  dma_read_addr13_to_bank16   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank16     =  read_request13_to_bank16    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank17
  wire dma_write_addr13_to_bank17      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr13_to_bank17       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank17   =  dma_write_addr13_to_bank17  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank17    =  write_request13_to_bank17   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank17    =  dma_read_addr13_to_bank17   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank17     =  read_request13_to_bank17    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank18
  wire dma_write_addr13_to_bank18      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr13_to_bank18       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank18   =  dma_write_addr13_to_bank18  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank18    =  write_request13_to_bank18   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank18    =  dma_read_addr13_to_bank18   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank18     =  read_request13_to_bank18    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank19
  wire dma_write_addr13_to_bank19      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr13_to_bank19       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank19   =  dma_write_addr13_to_bank19  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank19    =  write_request13_to_bank19   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank19    =  dma_read_addr13_to_bank19   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank19     =  read_request13_to_bank19    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank20
  wire dma_write_addr13_to_bank20      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr13_to_bank20       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank20   =  dma_write_addr13_to_bank20  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank20    =  write_request13_to_bank20   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank20    =  dma_read_addr13_to_bank20   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank20     =  read_request13_to_bank20    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank21
  wire dma_write_addr13_to_bank21      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr13_to_bank21       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank21   =  dma_write_addr13_to_bank21  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank21    =  write_request13_to_bank21   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank21    =  dma_read_addr13_to_bank21   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank21     =  read_request13_to_bank21    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank22
  wire dma_write_addr13_to_bank22      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr13_to_bank22       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank22   =  dma_write_addr13_to_bank22  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank22    =  write_request13_to_bank22   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank22    =  dma_read_addr13_to_bank22   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank22     =  read_request13_to_bank22    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank23
  wire dma_write_addr13_to_bank23      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr13_to_bank23       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank23   =  dma_write_addr13_to_bank23  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank23    =  write_request13_to_bank23   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank23    =  dma_read_addr13_to_bank23   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank23     =  read_request13_to_bank23    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank24
  wire dma_write_addr13_to_bank24      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr13_to_bank24       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank24   =  dma_write_addr13_to_bank24  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank24    =  write_request13_to_bank24   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank24    =  dma_read_addr13_to_bank24   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank24     =  read_request13_to_bank24    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank25
  wire dma_write_addr13_to_bank25      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr13_to_bank25       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank25   =  dma_write_addr13_to_bank25  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank25    =  write_request13_to_bank25   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank25    =  dma_read_addr13_to_bank25   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank25     =  read_request13_to_bank25    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank26
  wire dma_write_addr13_to_bank26      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr13_to_bank26       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank26   =  dma_write_addr13_to_bank26  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank26    =  write_request13_to_bank26   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank26    =  dma_read_addr13_to_bank26   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank26     =  read_request13_to_bank26    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank27
  wire dma_write_addr13_to_bank27      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr13_to_bank27       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank27   =  dma_write_addr13_to_bank27  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank27    =  write_request13_to_bank27   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank27    =  dma_read_addr13_to_bank27   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank27     =  read_request13_to_bank27    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank28
  wire dma_write_addr13_to_bank28      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr13_to_bank28       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank28   =  dma_write_addr13_to_bank28  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank28    =  write_request13_to_bank28   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank28    =  dma_read_addr13_to_bank28   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank28     =  read_request13_to_bank28    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank29
  wire dma_write_addr13_to_bank29      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr13_to_bank29       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank29   =  dma_write_addr13_to_bank29  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank29    =  write_request13_to_bank29   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank29    =  dma_read_addr13_to_bank29   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank29     =  read_request13_to_bank29    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank30
  wire dma_write_addr13_to_bank30      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr13_to_bank30       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank30   =  dma_write_addr13_to_bank30  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank30    =  write_request13_to_bank30   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank30    =  dma_read_addr13_to_bank30   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank30     =  read_request13_to_bank30    & memc__dma__read_ready13   ;                                         
  // DMA 13, bank31
  wire dma_write_addr13_to_bank31      =  (dma__memc__write_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr13_to_bank31       =  (dma__memc__read_address13[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank31   =  dma_write_addr13_to_bank31  & dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank31    =  write_request13_to_bank31   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank31    =  dma_read_addr13_to_bank31   & dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank31     =  read_request13_to_bank31    & memc__dma__read_ready13   ;                                         
  // DMA 14
  wire read_pause14     =  dma__memc__read_pause14   ;  
  // DMA 14, bank0
  wire dma_write_addr14_to_bank0      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr14_to_bank0       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank0   =  dma_write_addr14_to_bank0  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank0    =  write_request14_to_bank0   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank0    =  dma_read_addr14_to_bank0   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank0     =  read_request14_to_bank0    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank1
  wire dma_write_addr14_to_bank1      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr14_to_bank1       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank1   =  dma_write_addr14_to_bank1  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank1    =  write_request14_to_bank1   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank1    =  dma_read_addr14_to_bank1   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank1     =  read_request14_to_bank1    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank2
  wire dma_write_addr14_to_bank2      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr14_to_bank2       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank2   =  dma_write_addr14_to_bank2  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank2    =  write_request14_to_bank2   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank2    =  dma_read_addr14_to_bank2   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank2     =  read_request14_to_bank2    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank3
  wire dma_write_addr14_to_bank3      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr14_to_bank3       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank3   =  dma_write_addr14_to_bank3  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank3    =  write_request14_to_bank3   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank3    =  dma_read_addr14_to_bank3   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank3     =  read_request14_to_bank3    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank4
  wire dma_write_addr14_to_bank4      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr14_to_bank4       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank4   =  dma_write_addr14_to_bank4  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank4    =  write_request14_to_bank4   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank4    =  dma_read_addr14_to_bank4   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank4     =  read_request14_to_bank4    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank5
  wire dma_write_addr14_to_bank5      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr14_to_bank5       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank5   =  dma_write_addr14_to_bank5  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank5    =  write_request14_to_bank5   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank5    =  dma_read_addr14_to_bank5   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank5     =  read_request14_to_bank5    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank6
  wire dma_write_addr14_to_bank6      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr14_to_bank6       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank6   =  dma_write_addr14_to_bank6  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank6    =  write_request14_to_bank6   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank6    =  dma_read_addr14_to_bank6   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank6     =  read_request14_to_bank6    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank7
  wire dma_write_addr14_to_bank7      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr14_to_bank7       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank7   =  dma_write_addr14_to_bank7  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank7    =  write_request14_to_bank7   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank7    =  dma_read_addr14_to_bank7   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank7     =  read_request14_to_bank7    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank8
  wire dma_write_addr14_to_bank8      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr14_to_bank8       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank8   =  dma_write_addr14_to_bank8  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank8    =  write_request14_to_bank8   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank8    =  dma_read_addr14_to_bank8   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank8     =  read_request14_to_bank8    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank9
  wire dma_write_addr14_to_bank9      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr14_to_bank9       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank9   =  dma_write_addr14_to_bank9  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank9    =  write_request14_to_bank9   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank9    =  dma_read_addr14_to_bank9   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank9     =  read_request14_to_bank9    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank10
  wire dma_write_addr14_to_bank10      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr14_to_bank10       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank10   =  dma_write_addr14_to_bank10  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank10    =  write_request14_to_bank10   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank10    =  dma_read_addr14_to_bank10   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank10     =  read_request14_to_bank10    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank11
  wire dma_write_addr14_to_bank11      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr14_to_bank11       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank11   =  dma_write_addr14_to_bank11  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank11    =  write_request14_to_bank11   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank11    =  dma_read_addr14_to_bank11   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank11     =  read_request14_to_bank11    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank12
  wire dma_write_addr14_to_bank12      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr14_to_bank12       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank12   =  dma_write_addr14_to_bank12  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank12    =  write_request14_to_bank12   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank12    =  dma_read_addr14_to_bank12   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank12     =  read_request14_to_bank12    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank13
  wire dma_write_addr14_to_bank13      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr14_to_bank13       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank13   =  dma_write_addr14_to_bank13  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank13    =  write_request14_to_bank13   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank13    =  dma_read_addr14_to_bank13   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank13     =  read_request14_to_bank13    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank14
  wire dma_write_addr14_to_bank14      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr14_to_bank14       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank14   =  dma_write_addr14_to_bank14  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank14    =  write_request14_to_bank14   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank14    =  dma_read_addr14_to_bank14   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank14     =  read_request14_to_bank14    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank15
  wire dma_write_addr14_to_bank15      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr14_to_bank15       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank15   =  dma_write_addr14_to_bank15  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank15    =  write_request14_to_bank15   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank15    =  dma_read_addr14_to_bank15   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank15     =  read_request14_to_bank15    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank16
  wire dma_write_addr14_to_bank16      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr14_to_bank16       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank16   =  dma_write_addr14_to_bank16  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank16    =  write_request14_to_bank16   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank16    =  dma_read_addr14_to_bank16   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank16     =  read_request14_to_bank16    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank17
  wire dma_write_addr14_to_bank17      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr14_to_bank17       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank17   =  dma_write_addr14_to_bank17  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank17    =  write_request14_to_bank17   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank17    =  dma_read_addr14_to_bank17   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank17     =  read_request14_to_bank17    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank18
  wire dma_write_addr14_to_bank18      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr14_to_bank18       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank18   =  dma_write_addr14_to_bank18  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank18    =  write_request14_to_bank18   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank18    =  dma_read_addr14_to_bank18   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank18     =  read_request14_to_bank18    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank19
  wire dma_write_addr14_to_bank19      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr14_to_bank19       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank19   =  dma_write_addr14_to_bank19  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank19    =  write_request14_to_bank19   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank19    =  dma_read_addr14_to_bank19   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank19     =  read_request14_to_bank19    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank20
  wire dma_write_addr14_to_bank20      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr14_to_bank20       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank20   =  dma_write_addr14_to_bank20  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank20    =  write_request14_to_bank20   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank20    =  dma_read_addr14_to_bank20   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank20     =  read_request14_to_bank20    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank21
  wire dma_write_addr14_to_bank21      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr14_to_bank21       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank21   =  dma_write_addr14_to_bank21  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank21    =  write_request14_to_bank21   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank21    =  dma_read_addr14_to_bank21   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank21     =  read_request14_to_bank21    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank22
  wire dma_write_addr14_to_bank22      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr14_to_bank22       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank22   =  dma_write_addr14_to_bank22  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank22    =  write_request14_to_bank22   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank22    =  dma_read_addr14_to_bank22   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank22     =  read_request14_to_bank22    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank23
  wire dma_write_addr14_to_bank23      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr14_to_bank23       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank23   =  dma_write_addr14_to_bank23  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank23    =  write_request14_to_bank23   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank23    =  dma_read_addr14_to_bank23   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank23     =  read_request14_to_bank23    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank24
  wire dma_write_addr14_to_bank24      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr14_to_bank24       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank24   =  dma_write_addr14_to_bank24  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank24    =  write_request14_to_bank24   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank24    =  dma_read_addr14_to_bank24   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank24     =  read_request14_to_bank24    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank25
  wire dma_write_addr14_to_bank25      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr14_to_bank25       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank25   =  dma_write_addr14_to_bank25  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank25    =  write_request14_to_bank25   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank25    =  dma_read_addr14_to_bank25   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank25     =  read_request14_to_bank25    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank26
  wire dma_write_addr14_to_bank26      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr14_to_bank26       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank26   =  dma_write_addr14_to_bank26  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank26    =  write_request14_to_bank26   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank26    =  dma_read_addr14_to_bank26   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank26     =  read_request14_to_bank26    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank27
  wire dma_write_addr14_to_bank27      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr14_to_bank27       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank27   =  dma_write_addr14_to_bank27  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank27    =  write_request14_to_bank27   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank27    =  dma_read_addr14_to_bank27   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank27     =  read_request14_to_bank27    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank28
  wire dma_write_addr14_to_bank28      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr14_to_bank28       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank28   =  dma_write_addr14_to_bank28  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank28    =  write_request14_to_bank28   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank28    =  dma_read_addr14_to_bank28   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank28     =  read_request14_to_bank28    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank29
  wire dma_write_addr14_to_bank29      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr14_to_bank29       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank29   =  dma_write_addr14_to_bank29  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank29    =  write_request14_to_bank29   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank29    =  dma_read_addr14_to_bank29   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank29     =  read_request14_to_bank29    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank30
  wire dma_write_addr14_to_bank30      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr14_to_bank30       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank30   =  dma_write_addr14_to_bank30  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank30    =  write_request14_to_bank30   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank30    =  dma_read_addr14_to_bank30   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank30     =  read_request14_to_bank30    & memc__dma__read_ready14   ;                                         
  // DMA 14, bank31
  wire dma_write_addr14_to_bank31      =  (dma__memc__write_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr14_to_bank31       =  (dma__memc__read_address14[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank31   =  dma_write_addr14_to_bank31  & dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank31    =  write_request14_to_bank31   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank31    =  dma_read_addr14_to_bank31   & dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank31     =  read_request14_to_bank31    & memc__dma__read_ready14   ;                                         
  // DMA 15
  wire read_pause15     =  dma__memc__read_pause15   ;  
  // DMA 15, bank0
  wire dma_write_addr15_to_bank0      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr15_to_bank0       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank0   =  dma_write_addr15_to_bank0  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank0    =  write_request15_to_bank0   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank0    =  dma_read_addr15_to_bank0   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank0     =  read_request15_to_bank0    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank1
  wire dma_write_addr15_to_bank1      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr15_to_bank1       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank1   =  dma_write_addr15_to_bank1  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank1    =  write_request15_to_bank1   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank1    =  dma_read_addr15_to_bank1   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank1     =  read_request15_to_bank1    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank2
  wire dma_write_addr15_to_bank2      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr15_to_bank2       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank2   =  dma_write_addr15_to_bank2  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank2    =  write_request15_to_bank2   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank2    =  dma_read_addr15_to_bank2   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank2     =  read_request15_to_bank2    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank3
  wire dma_write_addr15_to_bank3      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr15_to_bank3       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank3   =  dma_write_addr15_to_bank3  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank3    =  write_request15_to_bank3   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank3    =  dma_read_addr15_to_bank3   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank3     =  read_request15_to_bank3    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank4
  wire dma_write_addr15_to_bank4      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr15_to_bank4       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank4   =  dma_write_addr15_to_bank4  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank4    =  write_request15_to_bank4   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank4    =  dma_read_addr15_to_bank4   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank4     =  read_request15_to_bank4    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank5
  wire dma_write_addr15_to_bank5      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr15_to_bank5       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank5   =  dma_write_addr15_to_bank5  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank5    =  write_request15_to_bank5   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank5    =  dma_read_addr15_to_bank5   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank5     =  read_request15_to_bank5    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank6
  wire dma_write_addr15_to_bank6      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr15_to_bank6       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank6   =  dma_write_addr15_to_bank6  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank6    =  write_request15_to_bank6   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank6    =  dma_read_addr15_to_bank6   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank6     =  read_request15_to_bank6    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank7
  wire dma_write_addr15_to_bank7      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr15_to_bank7       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank7   =  dma_write_addr15_to_bank7  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank7    =  write_request15_to_bank7   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank7    =  dma_read_addr15_to_bank7   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank7     =  read_request15_to_bank7    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank8
  wire dma_write_addr15_to_bank8      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr15_to_bank8       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank8   =  dma_write_addr15_to_bank8  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank8    =  write_request15_to_bank8   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank8    =  dma_read_addr15_to_bank8   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank8     =  read_request15_to_bank8    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank9
  wire dma_write_addr15_to_bank9      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr15_to_bank9       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank9   =  dma_write_addr15_to_bank9  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank9    =  write_request15_to_bank9   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank9    =  dma_read_addr15_to_bank9   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank9     =  read_request15_to_bank9    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank10
  wire dma_write_addr15_to_bank10      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr15_to_bank10       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank10   =  dma_write_addr15_to_bank10  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank10    =  write_request15_to_bank10   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank10    =  dma_read_addr15_to_bank10   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank10     =  read_request15_to_bank10    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank11
  wire dma_write_addr15_to_bank11      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr15_to_bank11       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank11   =  dma_write_addr15_to_bank11  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank11    =  write_request15_to_bank11   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank11    =  dma_read_addr15_to_bank11   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank11     =  read_request15_to_bank11    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank12
  wire dma_write_addr15_to_bank12      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr15_to_bank12       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank12   =  dma_write_addr15_to_bank12  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank12    =  write_request15_to_bank12   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank12    =  dma_read_addr15_to_bank12   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank12     =  read_request15_to_bank12    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank13
  wire dma_write_addr15_to_bank13      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr15_to_bank13       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank13   =  dma_write_addr15_to_bank13  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank13    =  write_request15_to_bank13   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank13    =  dma_read_addr15_to_bank13   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank13     =  read_request15_to_bank13    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank14
  wire dma_write_addr15_to_bank14      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr15_to_bank14       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank14   =  dma_write_addr15_to_bank14  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank14    =  write_request15_to_bank14   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank14    =  dma_read_addr15_to_bank14   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank14     =  read_request15_to_bank14    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank15
  wire dma_write_addr15_to_bank15      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr15_to_bank15       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank15   =  dma_write_addr15_to_bank15  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank15    =  write_request15_to_bank15   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank15    =  dma_read_addr15_to_bank15   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank15     =  read_request15_to_bank15    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank16
  wire dma_write_addr15_to_bank16      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr15_to_bank16       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank16   =  dma_write_addr15_to_bank16  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank16    =  write_request15_to_bank16   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank16    =  dma_read_addr15_to_bank16   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank16     =  read_request15_to_bank16    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank17
  wire dma_write_addr15_to_bank17      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr15_to_bank17       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank17   =  dma_write_addr15_to_bank17  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank17    =  write_request15_to_bank17   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank17    =  dma_read_addr15_to_bank17   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank17     =  read_request15_to_bank17    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank18
  wire dma_write_addr15_to_bank18      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr15_to_bank18       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank18   =  dma_write_addr15_to_bank18  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank18    =  write_request15_to_bank18   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank18    =  dma_read_addr15_to_bank18   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank18     =  read_request15_to_bank18    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank19
  wire dma_write_addr15_to_bank19      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr15_to_bank19       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank19   =  dma_write_addr15_to_bank19  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank19    =  write_request15_to_bank19   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank19    =  dma_read_addr15_to_bank19   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank19     =  read_request15_to_bank19    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank20
  wire dma_write_addr15_to_bank20      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr15_to_bank20       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank20   =  dma_write_addr15_to_bank20  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank20    =  write_request15_to_bank20   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank20    =  dma_read_addr15_to_bank20   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank20     =  read_request15_to_bank20    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank21
  wire dma_write_addr15_to_bank21      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr15_to_bank21       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank21   =  dma_write_addr15_to_bank21  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank21    =  write_request15_to_bank21   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank21    =  dma_read_addr15_to_bank21   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank21     =  read_request15_to_bank21    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank22
  wire dma_write_addr15_to_bank22      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr15_to_bank22       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank22   =  dma_write_addr15_to_bank22  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank22    =  write_request15_to_bank22   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank22    =  dma_read_addr15_to_bank22   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank22     =  read_request15_to_bank22    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank23
  wire dma_write_addr15_to_bank23      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr15_to_bank23       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank23   =  dma_write_addr15_to_bank23  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank23    =  write_request15_to_bank23   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank23    =  dma_read_addr15_to_bank23   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank23     =  read_request15_to_bank23    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank24
  wire dma_write_addr15_to_bank24      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr15_to_bank24       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank24   =  dma_write_addr15_to_bank24  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank24    =  write_request15_to_bank24   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank24    =  dma_read_addr15_to_bank24   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank24     =  read_request15_to_bank24    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank25
  wire dma_write_addr15_to_bank25      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr15_to_bank25       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank25   =  dma_write_addr15_to_bank25  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank25    =  write_request15_to_bank25   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank25    =  dma_read_addr15_to_bank25   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank25     =  read_request15_to_bank25    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank26
  wire dma_write_addr15_to_bank26      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr15_to_bank26       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank26   =  dma_write_addr15_to_bank26  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank26    =  write_request15_to_bank26   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank26    =  dma_read_addr15_to_bank26   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank26     =  read_request15_to_bank26    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank27
  wire dma_write_addr15_to_bank27      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr15_to_bank27       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank27   =  dma_write_addr15_to_bank27  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank27    =  write_request15_to_bank27   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank27    =  dma_read_addr15_to_bank27   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank27     =  read_request15_to_bank27    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank28
  wire dma_write_addr15_to_bank28      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr15_to_bank28       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank28   =  dma_write_addr15_to_bank28  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank28    =  write_request15_to_bank28   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank28    =  dma_read_addr15_to_bank28   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank28     =  read_request15_to_bank28    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank29
  wire dma_write_addr15_to_bank29      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr15_to_bank29       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank29   =  dma_write_addr15_to_bank29  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank29    =  write_request15_to_bank29   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank29    =  dma_read_addr15_to_bank29   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank29     =  read_request15_to_bank29    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank30
  wire dma_write_addr15_to_bank30      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr15_to_bank30       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank30   =  dma_write_addr15_to_bank30  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank30    =  write_request15_to_bank30   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank30    =  dma_read_addr15_to_bank30   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank30     =  read_request15_to_bank30    & memc__dma__read_ready15   ;                                         
  // DMA 15, bank31
  wire dma_write_addr15_to_bank31      =  (dma__memc__write_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr15_to_bank31       =  (dma__memc__read_address15[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank31   =  dma_write_addr15_to_bank31  & dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank31    =  write_request15_to_bank31   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank31    =  dma_read_addr15_to_bank31   & dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank31     =  read_request15_to_bank31    & memc__dma__read_ready15   ;                                         
  // DMA 16
  wire read_pause16     =  dma__memc__read_pause16   ;  
  // DMA 16, bank0
  wire dma_write_addr16_to_bank0      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr16_to_bank0       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank0   =  dma_write_addr16_to_bank0  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank0    =  write_request16_to_bank0   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank0    =  dma_read_addr16_to_bank0   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank0     =  read_request16_to_bank0    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank1
  wire dma_write_addr16_to_bank1      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr16_to_bank1       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank1   =  dma_write_addr16_to_bank1  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank1    =  write_request16_to_bank1   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank1    =  dma_read_addr16_to_bank1   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank1     =  read_request16_to_bank1    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank2
  wire dma_write_addr16_to_bank2      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr16_to_bank2       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank2   =  dma_write_addr16_to_bank2  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank2    =  write_request16_to_bank2   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank2    =  dma_read_addr16_to_bank2   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank2     =  read_request16_to_bank2    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank3
  wire dma_write_addr16_to_bank3      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr16_to_bank3       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank3   =  dma_write_addr16_to_bank3  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank3    =  write_request16_to_bank3   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank3    =  dma_read_addr16_to_bank3   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank3     =  read_request16_to_bank3    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank4
  wire dma_write_addr16_to_bank4      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr16_to_bank4       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank4   =  dma_write_addr16_to_bank4  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank4    =  write_request16_to_bank4   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank4    =  dma_read_addr16_to_bank4   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank4     =  read_request16_to_bank4    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank5
  wire dma_write_addr16_to_bank5      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr16_to_bank5       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank5   =  dma_write_addr16_to_bank5  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank5    =  write_request16_to_bank5   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank5    =  dma_read_addr16_to_bank5   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank5     =  read_request16_to_bank5    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank6
  wire dma_write_addr16_to_bank6      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr16_to_bank6       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank6   =  dma_write_addr16_to_bank6  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank6    =  write_request16_to_bank6   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank6    =  dma_read_addr16_to_bank6   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank6     =  read_request16_to_bank6    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank7
  wire dma_write_addr16_to_bank7      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr16_to_bank7       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank7   =  dma_write_addr16_to_bank7  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank7    =  write_request16_to_bank7   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank7    =  dma_read_addr16_to_bank7   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank7     =  read_request16_to_bank7    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank8
  wire dma_write_addr16_to_bank8      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr16_to_bank8       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank8   =  dma_write_addr16_to_bank8  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank8    =  write_request16_to_bank8   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank8    =  dma_read_addr16_to_bank8   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank8     =  read_request16_to_bank8    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank9
  wire dma_write_addr16_to_bank9      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr16_to_bank9       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank9   =  dma_write_addr16_to_bank9  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank9    =  write_request16_to_bank9   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank9    =  dma_read_addr16_to_bank9   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank9     =  read_request16_to_bank9    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank10
  wire dma_write_addr16_to_bank10      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr16_to_bank10       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank10   =  dma_write_addr16_to_bank10  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank10    =  write_request16_to_bank10   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank10    =  dma_read_addr16_to_bank10   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank10     =  read_request16_to_bank10    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank11
  wire dma_write_addr16_to_bank11      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr16_to_bank11       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank11   =  dma_write_addr16_to_bank11  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank11    =  write_request16_to_bank11   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank11    =  dma_read_addr16_to_bank11   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank11     =  read_request16_to_bank11    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank12
  wire dma_write_addr16_to_bank12      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr16_to_bank12       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank12   =  dma_write_addr16_to_bank12  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank12    =  write_request16_to_bank12   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank12    =  dma_read_addr16_to_bank12   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank12     =  read_request16_to_bank12    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank13
  wire dma_write_addr16_to_bank13      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr16_to_bank13       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank13   =  dma_write_addr16_to_bank13  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank13    =  write_request16_to_bank13   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank13    =  dma_read_addr16_to_bank13   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank13     =  read_request16_to_bank13    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank14
  wire dma_write_addr16_to_bank14      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr16_to_bank14       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank14   =  dma_write_addr16_to_bank14  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank14    =  write_request16_to_bank14   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank14    =  dma_read_addr16_to_bank14   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank14     =  read_request16_to_bank14    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank15
  wire dma_write_addr16_to_bank15      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr16_to_bank15       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank15   =  dma_write_addr16_to_bank15  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank15    =  write_request16_to_bank15   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank15    =  dma_read_addr16_to_bank15   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank15     =  read_request16_to_bank15    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank16
  wire dma_write_addr16_to_bank16      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr16_to_bank16       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank16   =  dma_write_addr16_to_bank16  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank16    =  write_request16_to_bank16   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank16    =  dma_read_addr16_to_bank16   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank16     =  read_request16_to_bank16    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank17
  wire dma_write_addr16_to_bank17      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr16_to_bank17       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank17   =  dma_write_addr16_to_bank17  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank17    =  write_request16_to_bank17   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank17    =  dma_read_addr16_to_bank17   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank17     =  read_request16_to_bank17    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank18
  wire dma_write_addr16_to_bank18      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr16_to_bank18       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank18   =  dma_write_addr16_to_bank18  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank18    =  write_request16_to_bank18   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank18    =  dma_read_addr16_to_bank18   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank18     =  read_request16_to_bank18    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank19
  wire dma_write_addr16_to_bank19      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr16_to_bank19       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank19   =  dma_write_addr16_to_bank19  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank19    =  write_request16_to_bank19   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank19    =  dma_read_addr16_to_bank19   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank19     =  read_request16_to_bank19    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank20
  wire dma_write_addr16_to_bank20      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr16_to_bank20       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank20   =  dma_write_addr16_to_bank20  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank20    =  write_request16_to_bank20   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank20    =  dma_read_addr16_to_bank20   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank20     =  read_request16_to_bank20    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank21
  wire dma_write_addr16_to_bank21      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr16_to_bank21       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank21   =  dma_write_addr16_to_bank21  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank21    =  write_request16_to_bank21   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank21    =  dma_read_addr16_to_bank21   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank21     =  read_request16_to_bank21    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank22
  wire dma_write_addr16_to_bank22      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr16_to_bank22       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank22   =  dma_write_addr16_to_bank22  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank22    =  write_request16_to_bank22   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank22    =  dma_read_addr16_to_bank22   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank22     =  read_request16_to_bank22    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank23
  wire dma_write_addr16_to_bank23      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr16_to_bank23       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank23   =  dma_write_addr16_to_bank23  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank23    =  write_request16_to_bank23   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank23    =  dma_read_addr16_to_bank23   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank23     =  read_request16_to_bank23    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank24
  wire dma_write_addr16_to_bank24      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr16_to_bank24       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank24   =  dma_write_addr16_to_bank24  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank24    =  write_request16_to_bank24   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank24    =  dma_read_addr16_to_bank24   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank24     =  read_request16_to_bank24    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank25
  wire dma_write_addr16_to_bank25      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr16_to_bank25       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank25   =  dma_write_addr16_to_bank25  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank25    =  write_request16_to_bank25   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank25    =  dma_read_addr16_to_bank25   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank25     =  read_request16_to_bank25    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank26
  wire dma_write_addr16_to_bank26      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr16_to_bank26       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank26   =  dma_write_addr16_to_bank26  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank26    =  write_request16_to_bank26   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank26    =  dma_read_addr16_to_bank26   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank26     =  read_request16_to_bank26    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank27
  wire dma_write_addr16_to_bank27      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr16_to_bank27       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank27   =  dma_write_addr16_to_bank27  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank27    =  write_request16_to_bank27   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank27    =  dma_read_addr16_to_bank27   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank27     =  read_request16_to_bank27    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank28
  wire dma_write_addr16_to_bank28      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr16_to_bank28       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank28   =  dma_write_addr16_to_bank28  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank28    =  write_request16_to_bank28   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank28    =  dma_read_addr16_to_bank28   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank28     =  read_request16_to_bank28    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank29
  wire dma_write_addr16_to_bank29      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr16_to_bank29       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank29   =  dma_write_addr16_to_bank29  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank29    =  write_request16_to_bank29   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank29    =  dma_read_addr16_to_bank29   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank29     =  read_request16_to_bank29    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank30
  wire dma_write_addr16_to_bank30      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr16_to_bank30       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank30   =  dma_write_addr16_to_bank30  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank30    =  write_request16_to_bank30   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank30    =  dma_read_addr16_to_bank30   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank30     =  read_request16_to_bank30    & memc__dma__read_ready16   ;                                         
  // DMA 16, bank31
  wire dma_write_addr16_to_bank31      =  (dma__memc__write_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr16_to_bank31       =  (dma__memc__read_address16[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank31   =  dma_write_addr16_to_bank31  & dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank31    =  write_request16_to_bank31   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank31    =  dma_read_addr16_to_bank31   & dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank31     =  read_request16_to_bank31    & memc__dma__read_ready16   ;                                         
  // DMA 17
  wire read_pause17     =  dma__memc__read_pause17   ;  
  // DMA 17, bank0
  wire dma_write_addr17_to_bank0      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr17_to_bank0       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank0   =  dma_write_addr17_to_bank0  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank0    =  write_request17_to_bank0   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank0    =  dma_read_addr17_to_bank0   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank0     =  read_request17_to_bank0    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank1
  wire dma_write_addr17_to_bank1      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr17_to_bank1       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank1   =  dma_write_addr17_to_bank1  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank1    =  write_request17_to_bank1   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank1    =  dma_read_addr17_to_bank1   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank1     =  read_request17_to_bank1    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank2
  wire dma_write_addr17_to_bank2      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr17_to_bank2       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank2   =  dma_write_addr17_to_bank2  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank2    =  write_request17_to_bank2   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank2    =  dma_read_addr17_to_bank2   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank2     =  read_request17_to_bank2    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank3
  wire dma_write_addr17_to_bank3      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr17_to_bank3       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank3   =  dma_write_addr17_to_bank3  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank3    =  write_request17_to_bank3   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank3    =  dma_read_addr17_to_bank3   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank3     =  read_request17_to_bank3    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank4
  wire dma_write_addr17_to_bank4      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr17_to_bank4       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank4   =  dma_write_addr17_to_bank4  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank4    =  write_request17_to_bank4   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank4    =  dma_read_addr17_to_bank4   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank4     =  read_request17_to_bank4    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank5
  wire dma_write_addr17_to_bank5      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr17_to_bank5       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank5   =  dma_write_addr17_to_bank5  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank5    =  write_request17_to_bank5   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank5    =  dma_read_addr17_to_bank5   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank5     =  read_request17_to_bank5    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank6
  wire dma_write_addr17_to_bank6      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr17_to_bank6       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank6   =  dma_write_addr17_to_bank6  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank6    =  write_request17_to_bank6   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank6    =  dma_read_addr17_to_bank6   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank6     =  read_request17_to_bank6    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank7
  wire dma_write_addr17_to_bank7      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr17_to_bank7       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank7   =  dma_write_addr17_to_bank7  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank7    =  write_request17_to_bank7   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank7    =  dma_read_addr17_to_bank7   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank7     =  read_request17_to_bank7    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank8
  wire dma_write_addr17_to_bank8      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr17_to_bank8       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank8   =  dma_write_addr17_to_bank8  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank8    =  write_request17_to_bank8   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank8    =  dma_read_addr17_to_bank8   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank8     =  read_request17_to_bank8    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank9
  wire dma_write_addr17_to_bank9      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr17_to_bank9       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank9   =  dma_write_addr17_to_bank9  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank9    =  write_request17_to_bank9   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank9    =  dma_read_addr17_to_bank9   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank9     =  read_request17_to_bank9    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank10
  wire dma_write_addr17_to_bank10      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr17_to_bank10       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank10   =  dma_write_addr17_to_bank10  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank10    =  write_request17_to_bank10   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank10    =  dma_read_addr17_to_bank10   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank10     =  read_request17_to_bank10    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank11
  wire dma_write_addr17_to_bank11      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr17_to_bank11       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank11   =  dma_write_addr17_to_bank11  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank11    =  write_request17_to_bank11   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank11    =  dma_read_addr17_to_bank11   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank11     =  read_request17_to_bank11    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank12
  wire dma_write_addr17_to_bank12      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr17_to_bank12       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank12   =  dma_write_addr17_to_bank12  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank12    =  write_request17_to_bank12   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank12    =  dma_read_addr17_to_bank12   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank12     =  read_request17_to_bank12    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank13
  wire dma_write_addr17_to_bank13      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr17_to_bank13       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank13   =  dma_write_addr17_to_bank13  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank13    =  write_request17_to_bank13   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank13    =  dma_read_addr17_to_bank13   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank13     =  read_request17_to_bank13    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank14
  wire dma_write_addr17_to_bank14      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr17_to_bank14       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank14   =  dma_write_addr17_to_bank14  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank14    =  write_request17_to_bank14   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank14    =  dma_read_addr17_to_bank14   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank14     =  read_request17_to_bank14    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank15
  wire dma_write_addr17_to_bank15      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr17_to_bank15       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank15   =  dma_write_addr17_to_bank15  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank15    =  write_request17_to_bank15   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank15    =  dma_read_addr17_to_bank15   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank15     =  read_request17_to_bank15    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank16
  wire dma_write_addr17_to_bank16      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr17_to_bank16       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank16   =  dma_write_addr17_to_bank16  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank16    =  write_request17_to_bank16   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank16    =  dma_read_addr17_to_bank16   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank16     =  read_request17_to_bank16    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank17
  wire dma_write_addr17_to_bank17      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr17_to_bank17       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank17   =  dma_write_addr17_to_bank17  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank17    =  write_request17_to_bank17   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank17    =  dma_read_addr17_to_bank17   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank17     =  read_request17_to_bank17    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank18
  wire dma_write_addr17_to_bank18      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr17_to_bank18       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank18   =  dma_write_addr17_to_bank18  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank18    =  write_request17_to_bank18   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank18    =  dma_read_addr17_to_bank18   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank18     =  read_request17_to_bank18    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank19
  wire dma_write_addr17_to_bank19      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr17_to_bank19       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank19   =  dma_write_addr17_to_bank19  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank19    =  write_request17_to_bank19   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank19    =  dma_read_addr17_to_bank19   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank19     =  read_request17_to_bank19    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank20
  wire dma_write_addr17_to_bank20      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr17_to_bank20       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank20   =  dma_write_addr17_to_bank20  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank20    =  write_request17_to_bank20   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank20    =  dma_read_addr17_to_bank20   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank20     =  read_request17_to_bank20    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank21
  wire dma_write_addr17_to_bank21      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr17_to_bank21       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank21   =  dma_write_addr17_to_bank21  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank21    =  write_request17_to_bank21   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank21    =  dma_read_addr17_to_bank21   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank21     =  read_request17_to_bank21    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank22
  wire dma_write_addr17_to_bank22      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr17_to_bank22       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank22   =  dma_write_addr17_to_bank22  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank22    =  write_request17_to_bank22   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank22    =  dma_read_addr17_to_bank22   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank22     =  read_request17_to_bank22    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank23
  wire dma_write_addr17_to_bank23      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr17_to_bank23       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank23   =  dma_write_addr17_to_bank23  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank23    =  write_request17_to_bank23   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank23    =  dma_read_addr17_to_bank23   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank23     =  read_request17_to_bank23    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank24
  wire dma_write_addr17_to_bank24      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr17_to_bank24       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank24   =  dma_write_addr17_to_bank24  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank24    =  write_request17_to_bank24   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank24    =  dma_read_addr17_to_bank24   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank24     =  read_request17_to_bank24    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank25
  wire dma_write_addr17_to_bank25      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr17_to_bank25       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank25   =  dma_write_addr17_to_bank25  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank25    =  write_request17_to_bank25   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank25    =  dma_read_addr17_to_bank25   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank25     =  read_request17_to_bank25    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank26
  wire dma_write_addr17_to_bank26      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr17_to_bank26       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank26   =  dma_write_addr17_to_bank26  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank26    =  write_request17_to_bank26   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank26    =  dma_read_addr17_to_bank26   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank26     =  read_request17_to_bank26    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank27
  wire dma_write_addr17_to_bank27      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr17_to_bank27       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank27   =  dma_write_addr17_to_bank27  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank27    =  write_request17_to_bank27   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank27    =  dma_read_addr17_to_bank27   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank27     =  read_request17_to_bank27    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank28
  wire dma_write_addr17_to_bank28      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr17_to_bank28       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank28   =  dma_write_addr17_to_bank28  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank28    =  write_request17_to_bank28   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank28    =  dma_read_addr17_to_bank28   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank28     =  read_request17_to_bank28    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank29
  wire dma_write_addr17_to_bank29      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr17_to_bank29       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank29   =  dma_write_addr17_to_bank29  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank29    =  write_request17_to_bank29   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank29    =  dma_read_addr17_to_bank29   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank29     =  read_request17_to_bank29    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank30
  wire dma_write_addr17_to_bank30      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr17_to_bank30       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank30   =  dma_write_addr17_to_bank30  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank30    =  write_request17_to_bank30   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank30    =  dma_read_addr17_to_bank30   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank30     =  read_request17_to_bank30    & memc__dma__read_ready17   ;                                         
  // DMA 17, bank31
  wire dma_write_addr17_to_bank31      =  (dma__memc__write_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr17_to_bank31       =  (dma__memc__read_address17[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank31   =  dma_write_addr17_to_bank31  & dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank31    =  write_request17_to_bank31   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank31    =  dma_read_addr17_to_bank31   & dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank31     =  read_request17_to_bank31    & memc__dma__read_ready17   ;                                         
  // DMA 18
  wire read_pause18     =  dma__memc__read_pause18   ;  
  // DMA 18, bank0
  wire dma_write_addr18_to_bank0      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr18_to_bank0       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank0   =  dma_write_addr18_to_bank0  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank0    =  write_request18_to_bank0   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank0    =  dma_read_addr18_to_bank0   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank0     =  read_request18_to_bank0    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank1
  wire dma_write_addr18_to_bank1      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr18_to_bank1       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank1   =  dma_write_addr18_to_bank1  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank1    =  write_request18_to_bank1   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank1    =  dma_read_addr18_to_bank1   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank1     =  read_request18_to_bank1    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank2
  wire dma_write_addr18_to_bank2      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr18_to_bank2       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank2   =  dma_write_addr18_to_bank2  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank2    =  write_request18_to_bank2   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank2    =  dma_read_addr18_to_bank2   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank2     =  read_request18_to_bank2    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank3
  wire dma_write_addr18_to_bank3      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr18_to_bank3       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank3   =  dma_write_addr18_to_bank3  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank3    =  write_request18_to_bank3   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank3    =  dma_read_addr18_to_bank3   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank3     =  read_request18_to_bank3    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank4
  wire dma_write_addr18_to_bank4      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr18_to_bank4       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank4   =  dma_write_addr18_to_bank4  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank4    =  write_request18_to_bank4   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank4    =  dma_read_addr18_to_bank4   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank4     =  read_request18_to_bank4    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank5
  wire dma_write_addr18_to_bank5      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr18_to_bank5       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank5   =  dma_write_addr18_to_bank5  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank5    =  write_request18_to_bank5   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank5    =  dma_read_addr18_to_bank5   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank5     =  read_request18_to_bank5    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank6
  wire dma_write_addr18_to_bank6      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr18_to_bank6       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank6   =  dma_write_addr18_to_bank6  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank6    =  write_request18_to_bank6   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank6    =  dma_read_addr18_to_bank6   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank6     =  read_request18_to_bank6    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank7
  wire dma_write_addr18_to_bank7      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr18_to_bank7       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank7   =  dma_write_addr18_to_bank7  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank7    =  write_request18_to_bank7   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank7    =  dma_read_addr18_to_bank7   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank7     =  read_request18_to_bank7    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank8
  wire dma_write_addr18_to_bank8      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr18_to_bank8       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank8   =  dma_write_addr18_to_bank8  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank8    =  write_request18_to_bank8   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank8    =  dma_read_addr18_to_bank8   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank8     =  read_request18_to_bank8    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank9
  wire dma_write_addr18_to_bank9      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr18_to_bank9       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank9   =  dma_write_addr18_to_bank9  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank9    =  write_request18_to_bank9   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank9    =  dma_read_addr18_to_bank9   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank9     =  read_request18_to_bank9    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank10
  wire dma_write_addr18_to_bank10      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr18_to_bank10       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank10   =  dma_write_addr18_to_bank10  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank10    =  write_request18_to_bank10   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank10    =  dma_read_addr18_to_bank10   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank10     =  read_request18_to_bank10    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank11
  wire dma_write_addr18_to_bank11      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr18_to_bank11       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank11   =  dma_write_addr18_to_bank11  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank11    =  write_request18_to_bank11   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank11    =  dma_read_addr18_to_bank11   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank11     =  read_request18_to_bank11    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank12
  wire dma_write_addr18_to_bank12      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr18_to_bank12       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank12   =  dma_write_addr18_to_bank12  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank12    =  write_request18_to_bank12   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank12    =  dma_read_addr18_to_bank12   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank12     =  read_request18_to_bank12    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank13
  wire dma_write_addr18_to_bank13      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr18_to_bank13       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank13   =  dma_write_addr18_to_bank13  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank13    =  write_request18_to_bank13   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank13    =  dma_read_addr18_to_bank13   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank13     =  read_request18_to_bank13    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank14
  wire dma_write_addr18_to_bank14      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr18_to_bank14       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank14   =  dma_write_addr18_to_bank14  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank14    =  write_request18_to_bank14   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank14    =  dma_read_addr18_to_bank14   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank14     =  read_request18_to_bank14    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank15
  wire dma_write_addr18_to_bank15      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr18_to_bank15       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank15   =  dma_write_addr18_to_bank15  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank15    =  write_request18_to_bank15   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank15    =  dma_read_addr18_to_bank15   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank15     =  read_request18_to_bank15    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank16
  wire dma_write_addr18_to_bank16      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr18_to_bank16       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank16   =  dma_write_addr18_to_bank16  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank16    =  write_request18_to_bank16   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank16    =  dma_read_addr18_to_bank16   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank16     =  read_request18_to_bank16    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank17
  wire dma_write_addr18_to_bank17      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr18_to_bank17       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank17   =  dma_write_addr18_to_bank17  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank17    =  write_request18_to_bank17   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank17    =  dma_read_addr18_to_bank17   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank17     =  read_request18_to_bank17    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank18
  wire dma_write_addr18_to_bank18      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr18_to_bank18       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank18   =  dma_write_addr18_to_bank18  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank18    =  write_request18_to_bank18   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank18    =  dma_read_addr18_to_bank18   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank18     =  read_request18_to_bank18    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank19
  wire dma_write_addr18_to_bank19      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr18_to_bank19       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank19   =  dma_write_addr18_to_bank19  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank19    =  write_request18_to_bank19   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank19    =  dma_read_addr18_to_bank19   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank19     =  read_request18_to_bank19    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank20
  wire dma_write_addr18_to_bank20      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr18_to_bank20       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank20   =  dma_write_addr18_to_bank20  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank20    =  write_request18_to_bank20   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank20    =  dma_read_addr18_to_bank20   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank20     =  read_request18_to_bank20    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank21
  wire dma_write_addr18_to_bank21      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr18_to_bank21       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank21   =  dma_write_addr18_to_bank21  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank21    =  write_request18_to_bank21   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank21    =  dma_read_addr18_to_bank21   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank21     =  read_request18_to_bank21    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank22
  wire dma_write_addr18_to_bank22      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr18_to_bank22       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank22   =  dma_write_addr18_to_bank22  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank22    =  write_request18_to_bank22   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank22    =  dma_read_addr18_to_bank22   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank22     =  read_request18_to_bank22    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank23
  wire dma_write_addr18_to_bank23      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr18_to_bank23       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank23   =  dma_write_addr18_to_bank23  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank23    =  write_request18_to_bank23   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank23    =  dma_read_addr18_to_bank23   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank23     =  read_request18_to_bank23    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank24
  wire dma_write_addr18_to_bank24      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr18_to_bank24       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank24   =  dma_write_addr18_to_bank24  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank24    =  write_request18_to_bank24   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank24    =  dma_read_addr18_to_bank24   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank24     =  read_request18_to_bank24    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank25
  wire dma_write_addr18_to_bank25      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr18_to_bank25       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank25   =  dma_write_addr18_to_bank25  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank25    =  write_request18_to_bank25   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank25    =  dma_read_addr18_to_bank25   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank25     =  read_request18_to_bank25    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank26
  wire dma_write_addr18_to_bank26      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr18_to_bank26       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank26   =  dma_write_addr18_to_bank26  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank26    =  write_request18_to_bank26   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank26    =  dma_read_addr18_to_bank26   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank26     =  read_request18_to_bank26    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank27
  wire dma_write_addr18_to_bank27      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr18_to_bank27       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank27   =  dma_write_addr18_to_bank27  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank27    =  write_request18_to_bank27   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank27    =  dma_read_addr18_to_bank27   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank27     =  read_request18_to_bank27    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank28
  wire dma_write_addr18_to_bank28      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr18_to_bank28       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank28   =  dma_write_addr18_to_bank28  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank28    =  write_request18_to_bank28   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank28    =  dma_read_addr18_to_bank28   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank28     =  read_request18_to_bank28    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank29
  wire dma_write_addr18_to_bank29      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr18_to_bank29       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank29   =  dma_write_addr18_to_bank29  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank29    =  write_request18_to_bank29   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank29    =  dma_read_addr18_to_bank29   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank29     =  read_request18_to_bank29    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank30
  wire dma_write_addr18_to_bank30      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr18_to_bank30       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank30   =  dma_write_addr18_to_bank30  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank30    =  write_request18_to_bank30   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank30    =  dma_read_addr18_to_bank30   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank30     =  read_request18_to_bank30    & memc__dma__read_ready18   ;                                         
  // DMA 18, bank31
  wire dma_write_addr18_to_bank31      =  (dma__memc__write_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr18_to_bank31       =  (dma__memc__read_address18[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank31   =  dma_write_addr18_to_bank31  & dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank31    =  write_request18_to_bank31   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank31    =  dma_read_addr18_to_bank31   & dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank31     =  read_request18_to_bank31    & memc__dma__read_ready18   ;                                         
  // DMA 19
  wire read_pause19     =  dma__memc__read_pause19   ;  
  // DMA 19, bank0
  wire dma_write_addr19_to_bank0      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr19_to_bank0       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank0   =  dma_write_addr19_to_bank0  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank0    =  write_request19_to_bank0   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank0    =  dma_read_addr19_to_bank0   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank0     =  read_request19_to_bank0    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank1
  wire dma_write_addr19_to_bank1      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr19_to_bank1       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank1   =  dma_write_addr19_to_bank1  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank1    =  write_request19_to_bank1   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank1    =  dma_read_addr19_to_bank1   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank1     =  read_request19_to_bank1    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank2
  wire dma_write_addr19_to_bank2      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr19_to_bank2       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank2   =  dma_write_addr19_to_bank2  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank2    =  write_request19_to_bank2   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank2    =  dma_read_addr19_to_bank2   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank2     =  read_request19_to_bank2    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank3
  wire dma_write_addr19_to_bank3      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr19_to_bank3       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank3   =  dma_write_addr19_to_bank3  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank3    =  write_request19_to_bank3   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank3    =  dma_read_addr19_to_bank3   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank3     =  read_request19_to_bank3    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank4
  wire dma_write_addr19_to_bank4      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr19_to_bank4       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank4   =  dma_write_addr19_to_bank4  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank4    =  write_request19_to_bank4   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank4    =  dma_read_addr19_to_bank4   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank4     =  read_request19_to_bank4    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank5
  wire dma_write_addr19_to_bank5      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr19_to_bank5       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank5   =  dma_write_addr19_to_bank5  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank5    =  write_request19_to_bank5   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank5    =  dma_read_addr19_to_bank5   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank5     =  read_request19_to_bank5    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank6
  wire dma_write_addr19_to_bank6      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr19_to_bank6       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank6   =  dma_write_addr19_to_bank6  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank6    =  write_request19_to_bank6   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank6    =  dma_read_addr19_to_bank6   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank6     =  read_request19_to_bank6    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank7
  wire dma_write_addr19_to_bank7      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr19_to_bank7       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank7   =  dma_write_addr19_to_bank7  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank7    =  write_request19_to_bank7   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank7    =  dma_read_addr19_to_bank7   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank7     =  read_request19_to_bank7    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank8
  wire dma_write_addr19_to_bank8      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr19_to_bank8       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank8   =  dma_write_addr19_to_bank8  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank8    =  write_request19_to_bank8   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank8    =  dma_read_addr19_to_bank8   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank8     =  read_request19_to_bank8    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank9
  wire dma_write_addr19_to_bank9      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr19_to_bank9       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank9   =  dma_write_addr19_to_bank9  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank9    =  write_request19_to_bank9   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank9    =  dma_read_addr19_to_bank9   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank9     =  read_request19_to_bank9    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank10
  wire dma_write_addr19_to_bank10      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr19_to_bank10       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank10   =  dma_write_addr19_to_bank10  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank10    =  write_request19_to_bank10   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank10    =  dma_read_addr19_to_bank10   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank10     =  read_request19_to_bank10    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank11
  wire dma_write_addr19_to_bank11      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr19_to_bank11       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank11   =  dma_write_addr19_to_bank11  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank11    =  write_request19_to_bank11   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank11    =  dma_read_addr19_to_bank11   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank11     =  read_request19_to_bank11    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank12
  wire dma_write_addr19_to_bank12      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr19_to_bank12       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank12   =  dma_write_addr19_to_bank12  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank12    =  write_request19_to_bank12   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank12    =  dma_read_addr19_to_bank12   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank12     =  read_request19_to_bank12    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank13
  wire dma_write_addr19_to_bank13      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr19_to_bank13       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank13   =  dma_write_addr19_to_bank13  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank13    =  write_request19_to_bank13   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank13    =  dma_read_addr19_to_bank13   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank13     =  read_request19_to_bank13    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank14
  wire dma_write_addr19_to_bank14      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr19_to_bank14       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank14   =  dma_write_addr19_to_bank14  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank14    =  write_request19_to_bank14   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank14    =  dma_read_addr19_to_bank14   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank14     =  read_request19_to_bank14    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank15
  wire dma_write_addr19_to_bank15      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr19_to_bank15       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank15   =  dma_write_addr19_to_bank15  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank15    =  write_request19_to_bank15   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank15    =  dma_read_addr19_to_bank15   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank15     =  read_request19_to_bank15    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank16
  wire dma_write_addr19_to_bank16      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr19_to_bank16       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank16   =  dma_write_addr19_to_bank16  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank16    =  write_request19_to_bank16   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank16    =  dma_read_addr19_to_bank16   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank16     =  read_request19_to_bank16    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank17
  wire dma_write_addr19_to_bank17      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr19_to_bank17       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank17   =  dma_write_addr19_to_bank17  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank17    =  write_request19_to_bank17   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank17    =  dma_read_addr19_to_bank17   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank17     =  read_request19_to_bank17    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank18
  wire dma_write_addr19_to_bank18      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr19_to_bank18       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank18   =  dma_write_addr19_to_bank18  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank18    =  write_request19_to_bank18   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank18    =  dma_read_addr19_to_bank18   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank18     =  read_request19_to_bank18    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank19
  wire dma_write_addr19_to_bank19      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr19_to_bank19       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank19   =  dma_write_addr19_to_bank19  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank19    =  write_request19_to_bank19   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank19    =  dma_read_addr19_to_bank19   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank19     =  read_request19_to_bank19    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank20
  wire dma_write_addr19_to_bank20      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr19_to_bank20       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank20   =  dma_write_addr19_to_bank20  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank20    =  write_request19_to_bank20   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank20    =  dma_read_addr19_to_bank20   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank20     =  read_request19_to_bank20    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank21
  wire dma_write_addr19_to_bank21      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr19_to_bank21       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank21   =  dma_write_addr19_to_bank21  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank21    =  write_request19_to_bank21   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank21    =  dma_read_addr19_to_bank21   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank21     =  read_request19_to_bank21    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank22
  wire dma_write_addr19_to_bank22      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr19_to_bank22       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank22   =  dma_write_addr19_to_bank22  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank22    =  write_request19_to_bank22   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank22    =  dma_read_addr19_to_bank22   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank22     =  read_request19_to_bank22    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank23
  wire dma_write_addr19_to_bank23      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr19_to_bank23       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank23   =  dma_write_addr19_to_bank23  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank23    =  write_request19_to_bank23   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank23    =  dma_read_addr19_to_bank23   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank23     =  read_request19_to_bank23    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank24
  wire dma_write_addr19_to_bank24      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr19_to_bank24       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank24   =  dma_write_addr19_to_bank24  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank24    =  write_request19_to_bank24   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank24    =  dma_read_addr19_to_bank24   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank24     =  read_request19_to_bank24    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank25
  wire dma_write_addr19_to_bank25      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr19_to_bank25       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank25   =  dma_write_addr19_to_bank25  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank25    =  write_request19_to_bank25   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank25    =  dma_read_addr19_to_bank25   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank25     =  read_request19_to_bank25    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank26
  wire dma_write_addr19_to_bank26      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr19_to_bank26       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank26   =  dma_write_addr19_to_bank26  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank26    =  write_request19_to_bank26   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank26    =  dma_read_addr19_to_bank26   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank26     =  read_request19_to_bank26    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank27
  wire dma_write_addr19_to_bank27      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr19_to_bank27       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank27   =  dma_write_addr19_to_bank27  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank27    =  write_request19_to_bank27   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank27    =  dma_read_addr19_to_bank27   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank27     =  read_request19_to_bank27    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank28
  wire dma_write_addr19_to_bank28      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr19_to_bank28       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank28   =  dma_write_addr19_to_bank28  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank28    =  write_request19_to_bank28   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank28    =  dma_read_addr19_to_bank28   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank28     =  read_request19_to_bank28    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank29
  wire dma_write_addr19_to_bank29      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr19_to_bank29       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank29   =  dma_write_addr19_to_bank29  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank29    =  write_request19_to_bank29   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank29    =  dma_read_addr19_to_bank29   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank29     =  read_request19_to_bank29    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank30
  wire dma_write_addr19_to_bank30      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr19_to_bank30       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank30   =  dma_write_addr19_to_bank30  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank30    =  write_request19_to_bank30   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank30    =  dma_read_addr19_to_bank30   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank30     =  read_request19_to_bank30    & memc__dma__read_ready19   ;                                         
  // DMA 19, bank31
  wire dma_write_addr19_to_bank31      =  (dma__memc__write_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr19_to_bank31       =  (dma__memc__read_address19[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank31   =  dma_write_addr19_to_bank31  & dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank31    =  write_request19_to_bank31   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank31    =  dma_read_addr19_to_bank31   & dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank31     =  read_request19_to_bank31    & memc__dma__read_ready19   ;                                         
  // DMA 20
  wire read_pause20     =  dma__memc__read_pause20   ;  
  // DMA 20, bank0
  wire dma_write_addr20_to_bank0      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr20_to_bank0       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank0   =  dma_write_addr20_to_bank0  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank0    =  write_request20_to_bank0   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank0    =  dma_read_addr20_to_bank0   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank0     =  read_request20_to_bank0    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank1
  wire dma_write_addr20_to_bank1      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr20_to_bank1       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank1   =  dma_write_addr20_to_bank1  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank1    =  write_request20_to_bank1   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank1    =  dma_read_addr20_to_bank1   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank1     =  read_request20_to_bank1    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank2
  wire dma_write_addr20_to_bank2      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr20_to_bank2       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank2   =  dma_write_addr20_to_bank2  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank2    =  write_request20_to_bank2   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank2    =  dma_read_addr20_to_bank2   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank2     =  read_request20_to_bank2    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank3
  wire dma_write_addr20_to_bank3      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr20_to_bank3       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank3   =  dma_write_addr20_to_bank3  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank3    =  write_request20_to_bank3   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank3    =  dma_read_addr20_to_bank3   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank3     =  read_request20_to_bank3    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank4
  wire dma_write_addr20_to_bank4      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr20_to_bank4       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank4   =  dma_write_addr20_to_bank4  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank4    =  write_request20_to_bank4   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank4    =  dma_read_addr20_to_bank4   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank4     =  read_request20_to_bank4    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank5
  wire dma_write_addr20_to_bank5      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr20_to_bank5       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank5   =  dma_write_addr20_to_bank5  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank5    =  write_request20_to_bank5   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank5    =  dma_read_addr20_to_bank5   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank5     =  read_request20_to_bank5    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank6
  wire dma_write_addr20_to_bank6      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr20_to_bank6       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank6   =  dma_write_addr20_to_bank6  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank6    =  write_request20_to_bank6   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank6    =  dma_read_addr20_to_bank6   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank6     =  read_request20_to_bank6    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank7
  wire dma_write_addr20_to_bank7      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr20_to_bank7       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank7   =  dma_write_addr20_to_bank7  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank7    =  write_request20_to_bank7   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank7    =  dma_read_addr20_to_bank7   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank7     =  read_request20_to_bank7    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank8
  wire dma_write_addr20_to_bank8      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr20_to_bank8       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank8   =  dma_write_addr20_to_bank8  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank8    =  write_request20_to_bank8   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank8    =  dma_read_addr20_to_bank8   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank8     =  read_request20_to_bank8    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank9
  wire dma_write_addr20_to_bank9      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr20_to_bank9       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank9   =  dma_write_addr20_to_bank9  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank9    =  write_request20_to_bank9   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank9    =  dma_read_addr20_to_bank9   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank9     =  read_request20_to_bank9    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank10
  wire dma_write_addr20_to_bank10      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr20_to_bank10       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank10   =  dma_write_addr20_to_bank10  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank10    =  write_request20_to_bank10   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank10    =  dma_read_addr20_to_bank10   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank10     =  read_request20_to_bank10    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank11
  wire dma_write_addr20_to_bank11      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr20_to_bank11       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank11   =  dma_write_addr20_to_bank11  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank11    =  write_request20_to_bank11   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank11    =  dma_read_addr20_to_bank11   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank11     =  read_request20_to_bank11    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank12
  wire dma_write_addr20_to_bank12      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr20_to_bank12       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank12   =  dma_write_addr20_to_bank12  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank12    =  write_request20_to_bank12   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank12    =  dma_read_addr20_to_bank12   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank12     =  read_request20_to_bank12    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank13
  wire dma_write_addr20_to_bank13      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr20_to_bank13       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank13   =  dma_write_addr20_to_bank13  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank13    =  write_request20_to_bank13   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank13    =  dma_read_addr20_to_bank13   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank13     =  read_request20_to_bank13    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank14
  wire dma_write_addr20_to_bank14      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr20_to_bank14       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank14   =  dma_write_addr20_to_bank14  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank14    =  write_request20_to_bank14   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank14    =  dma_read_addr20_to_bank14   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank14     =  read_request20_to_bank14    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank15
  wire dma_write_addr20_to_bank15      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr20_to_bank15       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank15   =  dma_write_addr20_to_bank15  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank15    =  write_request20_to_bank15   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank15    =  dma_read_addr20_to_bank15   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank15     =  read_request20_to_bank15    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank16
  wire dma_write_addr20_to_bank16      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr20_to_bank16       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank16   =  dma_write_addr20_to_bank16  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank16    =  write_request20_to_bank16   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank16    =  dma_read_addr20_to_bank16   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank16     =  read_request20_to_bank16    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank17
  wire dma_write_addr20_to_bank17      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr20_to_bank17       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank17   =  dma_write_addr20_to_bank17  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank17    =  write_request20_to_bank17   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank17    =  dma_read_addr20_to_bank17   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank17     =  read_request20_to_bank17    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank18
  wire dma_write_addr20_to_bank18      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr20_to_bank18       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank18   =  dma_write_addr20_to_bank18  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank18    =  write_request20_to_bank18   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank18    =  dma_read_addr20_to_bank18   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank18     =  read_request20_to_bank18    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank19
  wire dma_write_addr20_to_bank19      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr20_to_bank19       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank19   =  dma_write_addr20_to_bank19  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank19    =  write_request20_to_bank19   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank19    =  dma_read_addr20_to_bank19   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank19     =  read_request20_to_bank19    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank20
  wire dma_write_addr20_to_bank20      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr20_to_bank20       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank20   =  dma_write_addr20_to_bank20  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank20    =  write_request20_to_bank20   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank20    =  dma_read_addr20_to_bank20   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank20     =  read_request20_to_bank20    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank21
  wire dma_write_addr20_to_bank21      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr20_to_bank21       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank21   =  dma_write_addr20_to_bank21  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank21    =  write_request20_to_bank21   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank21    =  dma_read_addr20_to_bank21   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank21     =  read_request20_to_bank21    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank22
  wire dma_write_addr20_to_bank22      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr20_to_bank22       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank22   =  dma_write_addr20_to_bank22  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank22    =  write_request20_to_bank22   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank22    =  dma_read_addr20_to_bank22   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank22     =  read_request20_to_bank22    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank23
  wire dma_write_addr20_to_bank23      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr20_to_bank23       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank23   =  dma_write_addr20_to_bank23  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank23    =  write_request20_to_bank23   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank23    =  dma_read_addr20_to_bank23   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank23     =  read_request20_to_bank23    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank24
  wire dma_write_addr20_to_bank24      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr20_to_bank24       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank24   =  dma_write_addr20_to_bank24  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank24    =  write_request20_to_bank24   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank24    =  dma_read_addr20_to_bank24   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank24     =  read_request20_to_bank24    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank25
  wire dma_write_addr20_to_bank25      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr20_to_bank25       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank25   =  dma_write_addr20_to_bank25  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank25    =  write_request20_to_bank25   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank25    =  dma_read_addr20_to_bank25   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank25     =  read_request20_to_bank25    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank26
  wire dma_write_addr20_to_bank26      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr20_to_bank26       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank26   =  dma_write_addr20_to_bank26  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank26    =  write_request20_to_bank26   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank26    =  dma_read_addr20_to_bank26   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank26     =  read_request20_to_bank26    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank27
  wire dma_write_addr20_to_bank27      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr20_to_bank27       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank27   =  dma_write_addr20_to_bank27  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank27    =  write_request20_to_bank27   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank27    =  dma_read_addr20_to_bank27   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank27     =  read_request20_to_bank27    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank28
  wire dma_write_addr20_to_bank28      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr20_to_bank28       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank28   =  dma_write_addr20_to_bank28  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank28    =  write_request20_to_bank28   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank28    =  dma_read_addr20_to_bank28   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank28     =  read_request20_to_bank28    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank29
  wire dma_write_addr20_to_bank29      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr20_to_bank29       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank29   =  dma_write_addr20_to_bank29  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank29    =  write_request20_to_bank29   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank29    =  dma_read_addr20_to_bank29   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank29     =  read_request20_to_bank29    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank30
  wire dma_write_addr20_to_bank30      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr20_to_bank30       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank30   =  dma_write_addr20_to_bank30  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank30    =  write_request20_to_bank30   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank30    =  dma_read_addr20_to_bank30   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank30     =  read_request20_to_bank30    & memc__dma__read_ready20   ;                                         
  // DMA 20, bank31
  wire dma_write_addr20_to_bank31      =  (dma__memc__write_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr20_to_bank31       =  (dma__memc__read_address20[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank31   =  dma_write_addr20_to_bank31  & dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank31    =  write_request20_to_bank31   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank31    =  dma_read_addr20_to_bank31   & dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank31     =  read_request20_to_bank31    & memc__dma__read_ready20   ;                                         
  // DMA 21
  wire read_pause21     =  dma__memc__read_pause21   ;  
  // DMA 21, bank0
  wire dma_write_addr21_to_bank0      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr21_to_bank0       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank0   =  dma_write_addr21_to_bank0  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank0    =  write_request21_to_bank0   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank0    =  dma_read_addr21_to_bank0   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank0     =  read_request21_to_bank0    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank1
  wire dma_write_addr21_to_bank1      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr21_to_bank1       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank1   =  dma_write_addr21_to_bank1  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank1    =  write_request21_to_bank1   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank1    =  dma_read_addr21_to_bank1   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank1     =  read_request21_to_bank1    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank2
  wire dma_write_addr21_to_bank2      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr21_to_bank2       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank2   =  dma_write_addr21_to_bank2  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank2    =  write_request21_to_bank2   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank2    =  dma_read_addr21_to_bank2   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank2     =  read_request21_to_bank2    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank3
  wire dma_write_addr21_to_bank3      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr21_to_bank3       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank3   =  dma_write_addr21_to_bank3  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank3    =  write_request21_to_bank3   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank3    =  dma_read_addr21_to_bank3   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank3     =  read_request21_to_bank3    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank4
  wire dma_write_addr21_to_bank4      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr21_to_bank4       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank4   =  dma_write_addr21_to_bank4  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank4    =  write_request21_to_bank4   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank4    =  dma_read_addr21_to_bank4   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank4     =  read_request21_to_bank4    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank5
  wire dma_write_addr21_to_bank5      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr21_to_bank5       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank5   =  dma_write_addr21_to_bank5  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank5    =  write_request21_to_bank5   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank5    =  dma_read_addr21_to_bank5   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank5     =  read_request21_to_bank5    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank6
  wire dma_write_addr21_to_bank6      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr21_to_bank6       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank6   =  dma_write_addr21_to_bank6  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank6    =  write_request21_to_bank6   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank6    =  dma_read_addr21_to_bank6   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank6     =  read_request21_to_bank6    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank7
  wire dma_write_addr21_to_bank7      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr21_to_bank7       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank7   =  dma_write_addr21_to_bank7  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank7    =  write_request21_to_bank7   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank7    =  dma_read_addr21_to_bank7   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank7     =  read_request21_to_bank7    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank8
  wire dma_write_addr21_to_bank8      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr21_to_bank8       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank8   =  dma_write_addr21_to_bank8  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank8    =  write_request21_to_bank8   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank8    =  dma_read_addr21_to_bank8   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank8     =  read_request21_to_bank8    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank9
  wire dma_write_addr21_to_bank9      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr21_to_bank9       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank9   =  dma_write_addr21_to_bank9  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank9    =  write_request21_to_bank9   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank9    =  dma_read_addr21_to_bank9   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank9     =  read_request21_to_bank9    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank10
  wire dma_write_addr21_to_bank10      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr21_to_bank10       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank10   =  dma_write_addr21_to_bank10  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank10    =  write_request21_to_bank10   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank10    =  dma_read_addr21_to_bank10   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank10     =  read_request21_to_bank10    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank11
  wire dma_write_addr21_to_bank11      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr21_to_bank11       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank11   =  dma_write_addr21_to_bank11  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank11    =  write_request21_to_bank11   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank11    =  dma_read_addr21_to_bank11   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank11     =  read_request21_to_bank11    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank12
  wire dma_write_addr21_to_bank12      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr21_to_bank12       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank12   =  dma_write_addr21_to_bank12  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank12    =  write_request21_to_bank12   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank12    =  dma_read_addr21_to_bank12   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank12     =  read_request21_to_bank12    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank13
  wire dma_write_addr21_to_bank13      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr21_to_bank13       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank13   =  dma_write_addr21_to_bank13  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank13    =  write_request21_to_bank13   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank13    =  dma_read_addr21_to_bank13   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank13     =  read_request21_to_bank13    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank14
  wire dma_write_addr21_to_bank14      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr21_to_bank14       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank14   =  dma_write_addr21_to_bank14  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank14    =  write_request21_to_bank14   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank14    =  dma_read_addr21_to_bank14   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank14     =  read_request21_to_bank14    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank15
  wire dma_write_addr21_to_bank15      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr21_to_bank15       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank15   =  dma_write_addr21_to_bank15  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank15    =  write_request21_to_bank15   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank15    =  dma_read_addr21_to_bank15   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank15     =  read_request21_to_bank15    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank16
  wire dma_write_addr21_to_bank16      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr21_to_bank16       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank16   =  dma_write_addr21_to_bank16  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank16    =  write_request21_to_bank16   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank16    =  dma_read_addr21_to_bank16   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank16     =  read_request21_to_bank16    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank17
  wire dma_write_addr21_to_bank17      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr21_to_bank17       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank17   =  dma_write_addr21_to_bank17  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank17    =  write_request21_to_bank17   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank17    =  dma_read_addr21_to_bank17   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank17     =  read_request21_to_bank17    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank18
  wire dma_write_addr21_to_bank18      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr21_to_bank18       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank18   =  dma_write_addr21_to_bank18  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank18    =  write_request21_to_bank18   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank18    =  dma_read_addr21_to_bank18   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank18     =  read_request21_to_bank18    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank19
  wire dma_write_addr21_to_bank19      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr21_to_bank19       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank19   =  dma_write_addr21_to_bank19  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank19    =  write_request21_to_bank19   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank19    =  dma_read_addr21_to_bank19   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank19     =  read_request21_to_bank19    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank20
  wire dma_write_addr21_to_bank20      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr21_to_bank20       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank20   =  dma_write_addr21_to_bank20  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank20    =  write_request21_to_bank20   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank20    =  dma_read_addr21_to_bank20   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank20     =  read_request21_to_bank20    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank21
  wire dma_write_addr21_to_bank21      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr21_to_bank21       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank21   =  dma_write_addr21_to_bank21  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank21    =  write_request21_to_bank21   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank21    =  dma_read_addr21_to_bank21   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank21     =  read_request21_to_bank21    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank22
  wire dma_write_addr21_to_bank22      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr21_to_bank22       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank22   =  dma_write_addr21_to_bank22  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank22    =  write_request21_to_bank22   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank22    =  dma_read_addr21_to_bank22   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank22     =  read_request21_to_bank22    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank23
  wire dma_write_addr21_to_bank23      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr21_to_bank23       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank23   =  dma_write_addr21_to_bank23  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank23    =  write_request21_to_bank23   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank23    =  dma_read_addr21_to_bank23   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank23     =  read_request21_to_bank23    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank24
  wire dma_write_addr21_to_bank24      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr21_to_bank24       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank24   =  dma_write_addr21_to_bank24  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank24    =  write_request21_to_bank24   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank24    =  dma_read_addr21_to_bank24   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank24     =  read_request21_to_bank24    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank25
  wire dma_write_addr21_to_bank25      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr21_to_bank25       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank25   =  dma_write_addr21_to_bank25  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank25    =  write_request21_to_bank25   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank25    =  dma_read_addr21_to_bank25   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank25     =  read_request21_to_bank25    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank26
  wire dma_write_addr21_to_bank26      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr21_to_bank26       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank26   =  dma_write_addr21_to_bank26  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank26    =  write_request21_to_bank26   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank26    =  dma_read_addr21_to_bank26   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank26     =  read_request21_to_bank26    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank27
  wire dma_write_addr21_to_bank27      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr21_to_bank27       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank27   =  dma_write_addr21_to_bank27  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank27    =  write_request21_to_bank27   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank27    =  dma_read_addr21_to_bank27   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank27     =  read_request21_to_bank27    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank28
  wire dma_write_addr21_to_bank28      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr21_to_bank28       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank28   =  dma_write_addr21_to_bank28  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank28    =  write_request21_to_bank28   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank28    =  dma_read_addr21_to_bank28   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank28     =  read_request21_to_bank28    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank29
  wire dma_write_addr21_to_bank29      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr21_to_bank29       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank29   =  dma_write_addr21_to_bank29  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank29    =  write_request21_to_bank29   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank29    =  dma_read_addr21_to_bank29   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank29     =  read_request21_to_bank29    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank30
  wire dma_write_addr21_to_bank30      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr21_to_bank30       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank30   =  dma_write_addr21_to_bank30  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank30    =  write_request21_to_bank30   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank30    =  dma_read_addr21_to_bank30   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank30     =  read_request21_to_bank30    & memc__dma__read_ready21   ;                                         
  // DMA 21, bank31
  wire dma_write_addr21_to_bank31      =  (dma__memc__write_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr21_to_bank31       =  (dma__memc__read_address21[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank31   =  dma_write_addr21_to_bank31  & dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank31    =  write_request21_to_bank31   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank31    =  dma_read_addr21_to_bank31   & dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank31     =  read_request21_to_bank31    & memc__dma__read_ready21   ;                                         
  // DMA 22
  wire read_pause22     =  dma__memc__read_pause22   ;  
  // DMA 22, bank0
  wire dma_write_addr22_to_bank0      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr22_to_bank0       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank0   =  dma_write_addr22_to_bank0  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank0    =  write_request22_to_bank0   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank0    =  dma_read_addr22_to_bank0   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank0     =  read_request22_to_bank0    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank1
  wire dma_write_addr22_to_bank1      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr22_to_bank1       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank1   =  dma_write_addr22_to_bank1  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank1    =  write_request22_to_bank1   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank1    =  dma_read_addr22_to_bank1   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank1     =  read_request22_to_bank1    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank2
  wire dma_write_addr22_to_bank2      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr22_to_bank2       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank2   =  dma_write_addr22_to_bank2  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank2    =  write_request22_to_bank2   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank2    =  dma_read_addr22_to_bank2   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank2     =  read_request22_to_bank2    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank3
  wire dma_write_addr22_to_bank3      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr22_to_bank3       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank3   =  dma_write_addr22_to_bank3  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank3    =  write_request22_to_bank3   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank3    =  dma_read_addr22_to_bank3   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank3     =  read_request22_to_bank3    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank4
  wire dma_write_addr22_to_bank4      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr22_to_bank4       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank4   =  dma_write_addr22_to_bank4  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank4    =  write_request22_to_bank4   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank4    =  dma_read_addr22_to_bank4   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank4     =  read_request22_to_bank4    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank5
  wire dma_write_addr22_to_bank5      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr22_to_bank5       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank5   =  dma_write_addr22_to_bank5  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank5    =  write_request22_to_bank5   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank5    =  dma_read_addr22_to_bank5   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank5     =  read_request22_to_bank5    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank6
  wire dma_write_addr22_to_bank6      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr22_to_bank6       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank6   =  dma_write_addr22_to_bank6  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank6    =  write_request22_to_bank6   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank6    =  dma_read_addr22_to_bank6   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank6     =  read_request22_to_bank6    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank7
  wire dma_write_addr22_to_bank7      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr22_to_bank7       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank7   =  dma_write_addr22_to_bank7  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank7    =  write_request22_to_bank7   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank7    =  dma_read_addr22_to_bank7   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank7     =  read_request22_to_bank7    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank8
  wire dma_write_addr22_to_bank8      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr22_to_bank8       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank8   =  dma_write_addr22_to_bank8  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank8    =  write_request22_to_bank8   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank8    =  dma_read_addr22_to_bank8   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank8     =  read_request22_to_bank8    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank9
  wire dma_write_addr22_to_bank9      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr22_to_bank9       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank9   =  dma_write_addr22_to_bank9  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank9    =  write_request22_to_bank9   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank9    =  dma_read_addr22_to_bank9   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank9     =  read_request22_to_bank9    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank10
  wire dma_write_addr22_to_bank10      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr22_to_bank10       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank10   =  dma_write_addr22_to_bank10  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank10    =  write_request22_to_bank10   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank10    =  dma_read_addr22_to_bank10   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank10     =  read_request22_to_bank10    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank11
  wire dma_write_addr22_to_bank11      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr22_to_bank11       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank11   =  dma_write_addr22_to_bank11  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank11    =  write_request22_to_bank11   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank11    =  dma_read_addr22_to_bank11   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank11     =  read_request22_to_bank11    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank12
  wire dma_write_addr22_to_bank12      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr22_to_bank12       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank12   =  dma_write_addr22_to_bank12  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank12    =  write_request22_to_bank12   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank12    =  dma_read_addr22_to_bank12   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank12     =  read_request22_to_bank12    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank13
  wire dma_write_addr22_to_bank13      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr22_to_bank13       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank13   =  dma_write_addr22_to_bank13  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank13    =  write_request22_to_bank13   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank13    =  dma_read_addr22_to_bank13   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank13     =  read_request22_to_bank13    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank14
  wire dma_write_addr22_to_bank14      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr22_to_bank14       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank14   =  dma_write_addr22_to_bank14  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank14    =  write_request22_to_bank14   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank14    =  dma_read_addr22_to_bank14   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank14     =  read_request22_to_bank14    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank15
  wire dma_write_addr22_to_bank15      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr22_to_bank15       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank15   =  dma_write_addr22_to_bank15  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank15    =  write_request22_to_bank15   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank15    =  dma_read_addr22_to_bank15   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank15     =  read_request22_to_bank15    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank16
  wire dma_write_addr22_to_bank16      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr22_to_bank16       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank16   =  dma_write_addr22_to_bank16  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank16    =  write_request22_to_bank16   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank16    =  dma_read_addr22_to_bank16   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank16     =  read_request22_to_bank16    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank17
  wire dma_write_addr22_to_bank17      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr22_to_bank17       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank17   =  dma_write_addr22_to_bank17  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank17    =  write_request22_to_bank17   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank17    =  dma_read_addr22_to_bank17   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank17     =  read_request22_to_bank17    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank18
  wire dma_write_addr22_to_bank18      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr22_to_bank18       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank18   =  dma_write_addr22_to_bank18  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank18    =  write_request22_to_bank18   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank18    =  dma_read_addr22_to_bank18   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank18     =  read_request22_to_bank18    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank19
  wire dma_write_addr22_to_bank19      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr22_to_bank19       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank19   =  dma_write_addr22_to_bank19  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank19    =  write_request22_to_bank19   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank19    =  dma_read_addr22_to_bank19   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank19     =  read_request22_to_bank19    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank20
  wire dma_write_addr22_to_bank20      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr22_to_bank20       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank20   =  dma_write_addr22_to_bank20  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank20    =  write_request22_to_bank20   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank20    =  dma_read_addr22_to_bank20   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank20     =  read_request22_to_bank20    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank21
  wire dma_write_addr22_to_bank21      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr22_to_bank21       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank21   =  dma_write_addr22_to_bank21  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank21    =  write_request22_to_bank21   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank21    =  dma_read_addr22_to_bank21   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank21     =  read_request22_to_bank21    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank22
  wire dma_write_addr22_to_bank22      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr22_to_bank22       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank22   =  dma_write_addr22_to_bank22  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank22    =  write_request22_to_bank22   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank22    =  dma_read_addr22_to_bank22   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank22     =  read_request22_to_bank22    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank23
  wire dma_write_addr22_to_bank23      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr22_to_bank23       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank23   =  dma_write_addr22_to_bank23  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank23    =  write_request22_to_bank23   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank23    =  dma_read_addr22_to_bank23   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank23     =  read_request22_to_bank23    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank24
  wire dma_write_addr22_to_bank24      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr22_to_bank24       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank24   =  dma_write_addr22_to_bank24  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank24    =  write_request22_to_bank24   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank24    =  dma_read_addr22_to_bank24   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank24     =  read_request22_to_bank24    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank25
  wire dma_write_addr22_to_bank25      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr22_to_bank25       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank25   =  dma_write_addr22_to_bank25  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank25    =  write_request22_to_bank25   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank25    =  dma_read_addr22_to_bank25   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank25     =  read_request22_to_bank25    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank26
  wire dma_write_addr22_to_bank26      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr22_to_bank26       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank26   =  dma_write_addr22_to_bank26  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank26    =  write_request22_to_bank26   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank26    =  dma_read_addr22_to_bank26   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank26     =  read_request22_to_bank26    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank27
  wire dma_write_addr22_to_bank27      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr22_to_bank27       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank27   =  dma_write_addr22_to_bank27  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank27    =  write_request22_to_bank27   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank27    =  dma_read_addr22_to_bank27   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank27     =  read_request22_to_bank27    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank28
  wire dma_write_addr22_to_bank28      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr22_to_bank28       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank28   =  dma_write_addr22_to_bank28  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank28    =  write_request22_to_bank28   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank28    =  dma_read_addr22_to_bank28   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank28     =  read_request22_to_bank28    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank29
  wire dma_write_addr22_to_bank29      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr22_to_bank29       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank29   =  dma_write_addr22_to_bank29  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank29    =  write_request22_to_bank29   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank29    =  dma_read_addr22_to_bank29   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank29     =  read_request22_to_bank29    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank30
  wire dma_write_addr22_to_bank30      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr22_to_bank30       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank30   =  dma_write_addr22_to_bank30  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank30    =  write_request22_to_bank30   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank30    =  dma_read_addr22_to_bank30   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank30     =  read_request22_to_bank30    & memc__dma__read_ready22   ;                                         
  // DMA 22, bank31
  wire dma_write_addr22_to_bank31      =  (dma__memc__write_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr22_to_bank31       =  (dma__memc__read_address22[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank31   =  dma_write_addr22_to_bank31  & dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank31    =  write_request22_to_bank31   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank31    =  dma_read_addr22_to_bank31   & dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank31     =  read_request22_to_bank31    & memc__dma__read_ready22   ;                                         
  // DMA 23
  wire read_pause23     =  dma__memc__read_pause23   ;  
  // DMA 23, bank0
  wire dma_write_addr23_to_bank0      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr23_to_bank0       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank0   =  dma_write_addr23_to_bank0  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank0    =  write_request23_to_bank0   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank0    =  dma_read_addr23_to_bank0   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank0     =  read_request23_to_bank0    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank1
  wire dma_write_addr23_to_bank1      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr23_to_bank1       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank1   =  dma_write_addr23_to_bank1  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank1    =  write_request23_to_bank1   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank1    =  dma_read_addr23_to_bank1   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank1     =  read_request23_to_bank1    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank2
  wire dma_write_addr23_to_bank2      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr23_to_bank2       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank2   =  dma_write_addr23_to_bank2  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank2    =  write_request23_to_bank2   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank2    =  dma_read_addr23_to_bank2   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank2     =  read_request23_to_bank2    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank3
  wire dma_write_addr23_to_bank3      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr23_to_bank3       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank3   =  dma_write_addr23_to_bank3  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank3    =  write_request23_to_bank3   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank3    =  dma_read_addr23_to_bank3   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank3     =  read_request23_to_bank3    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank4
  wire dma_write_addr23_to_bank4      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr23_to_bank4       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank4   =  dma_write_addr23_to_bank4  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank4    =  write_request23_to_bank4   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank4    =  dma_read_addr23_to_bank4   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank4     =  read_request23_to_bank4    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank5
  wire dma_write_addr23_to_bank5      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr23_to_bank5       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank5   =  dma_write_addr23_to_bank5  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank5    =  write_request23_to_bank5   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank5    =  dma_read_addr23_to_bank5   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank5     =  read_request23_to_bank5    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank6
  wire dma_write_addr23_to_bank6      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr23_to_bank6       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank6   =  dma_write_addr23_to_bank6  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank6    =  write_request23_to_bank6   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank6    =  dma_read_addr23_to_bank6   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank6     =  read_request23_to_bank6    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank7
  wire dma_write_addr23_to_bank7      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr23_to_bank7       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank7   =  dma_write_addr23_to_bank7  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank7    =  write_request23_to_bank7   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank7    =  dma_read_addr23_to_bank7   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank7     =  read_request23_to_bank7    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank8
  wire dma_write_addr23_to_bank8      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr23_to_bank8       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank8   =  dma_write_addr23_to_bank8  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank8    =  write_request23_to_bank8   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank8    =  dma_read_addr23_to_bank8   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank8     =  read_request23_to_bank8    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank9
  wire dma_write_addr23_to_bank9      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr23_to_bank9       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank9   =  dma_write_addr23_to_bank9  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank9    =  write_request23_to_bank9   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank9    =  dma_read_addr23_to_bank9   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank9     =  read_request23_to_bank9    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank10
  wire dma_write_addr23_to_bank10      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr23_to_bank10       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank10   =  dma_write_addr23_to_bank10  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank10    =  write_request23_to_bank10   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank10    =  dma_read_addr23_to_bank10   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank10     =  read_request23_to_bank10    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank11
  wire dma_write_addr23_to_bank11      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr23_to_bank11       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank11   =  dma_write_addr23_to_bank11  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank11    =  write_request23_to_bank11   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank11    =  dma_read_addr23_to_bank11   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank11     =  read_request23_to_bank11    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank12
  wire dma_write_addr23_to_bank12      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr23_to_bank12       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank12   =  dma_write_addr23_to_bank12  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank12    =  write_request23_to_bank12   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank12    =  dma_read_addr23_to_bank12   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank12     =  read_request23_to_bank12    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank13
  wire dma_write_addr23_to_bank13      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr23_to_bank13       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank13   =  dma_write_addr23_to_bank13  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank13    =  write_request23_to_bank13   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank13    =  dma_read_addr23_to_bank13   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank13     =  read_request23_to_bank13    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank14
  wire dma_write_addr23_to_bank14      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr23_to_bank14       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank14   =  dma_write_addr23_to_bank14  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank14    =  write_request23_to_bank14   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank14    =  dma_read_addr23_to_bank14   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank14     =  read_request23_to_bank14    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank15
  wire dma_write_addr23_to_bank15      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr23_to_bank15       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank15   =  dma_write_addr23_to_bank15  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank15    =  write_request23_to_bank15   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank15    =  dma_read_addr23_to_bank15   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank15     =  read_request23_to_bank15    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank16
  wire dma_write_addr23_to_bank16      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr23_to_bank16       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank16   =  dma_write_addr23_to_bank16  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank16    =  write_request23_to_bank16   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank16    =  dma_read_addr23_to_bank16   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank16     =  read_request23_to_bank16    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank17
  wire dma_write_addr23_to_bank17      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr23_to_bank17       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank17   =  dma_write_addr23_to_bank17  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank17    =  write_request23_to_bank17   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank17    =  dma_read_addr23_to_bank17   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank17     =  read_request23_to_bank17    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank18
  wire dma_write_addr23_to_bank18      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr23_to_bank18       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank18   =  dma_write_addr23_to_bank18  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank18    =  write_request23_to_bank18   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank18    =  dma_read_addr23_to_bank18   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank18     =  read_request23_to_bank18    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank19
  wire dma_write_addr23_to_bank19      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr23_to_bank19       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank19   =  dma_write_addr23_to_bank19  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank19    =  write_request23_to_bank19   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank19    =  dma_read_addr23_to_bank19   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank19     =  read_request23_to_bank19    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank20
  wire dma_write_addr23_to_bank20      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr23_to_bank20       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank20   =  dma_write_addr23_to_bank20  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank20    =  write_request23_to_bank20   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank20    =  dma_read_addr23_to_bank20   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank20     =  read_request23_to_bank20    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank21
  wire dma_write_addr23_to_bank21      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr23_to_bank21       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank21   =  dma_write_addr23_to_bank21  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank21    =  write_request23_to_bank21   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank21    =  dma_read_addr23_to_bank21   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank21     =  read_request23_to_bank21    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank22
  wire dma_write_addr23_to_bank22      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr23_to_bank22       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank22   =  dma_write_addr23_to_bank22  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank22    =  write_request23_to_bank22   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank22    =  dma_read_addr23_to_bank22   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank22     =  read_request23_to_bank22    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank23
  wire dma_write_addr23_to_bank23      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr23_to_bank23       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank23   =  dma_write_addr23_to_bank23  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank23    =  write_request23_to_bank23   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank23    =  dma_read_addr23_to_bank23   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank23     =  read_request23_to_bank23    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank24
  wire dma_write_addr23_to_bank24      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr23_to_bank24       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank24   =  dma_write_addr23_to_bank24  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank24    =  write_request23_to_bank24   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank24    =  dma_read_addr23_to_bank24   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank24     =  read_request23_to_bank24    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank25
  wire dma_write_addr23_to_bank25      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr23_to_bank25       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank25   =  dma_write_addr23_to_bank25  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank25    =  write_request23_to_bank25   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank25    =  dma_read_addr23_to_bank25   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank25     =  read_request23_to_bank25    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank26
  wire dma_write_addr23_to_bank26      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr23_to_bank26       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank26   =  dma_write_addr23_to_bank26  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank26    =  write_request23_to_bank26   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank26    =  dma_read_addr23_to_bank26   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank26     =  read_request23_to_bank26    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank27
  wire dma_write_addr23_to_bank27      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr23_to_bank27       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank27   =  dma_write_addr23_to_bank27  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank27    =  write_request23_to_bank27   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank27    =  dma_read_addr23_to_bank27   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank27     =  read_request23_to_bank27    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank28
  wire dma_write_addr23_to_bank28      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr23_to_bank28       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank28   =  dma_write_addr23_to_bank28  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank28    =  write_request23_to_bank28   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank28    =  dma_read_addr23_to_bank28   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank28     =  read_request23_to_bank28    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank29
  wire dma_write_addr23_to_bank29      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr23_to_bank29       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank29   =  dma_write_addr23_to_bank29  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank29    =  write_request23_to_bank29   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank29    =  dma_read_addr23_to_bank29   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank29     =  read_request23_to_bank29    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank30
  wire dma_write_addr23_to_bank30      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr23_to_bank30       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank30   =  dma_write_addr23_to_bank30  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank30    =  write_request23_to_bank30   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank30    =  dma_read_addr23_to_bank30   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank30     =  read_request23_to_bank30    & memc__dma__read_ready23   ;                                         
  // DMA 23, bank31
  wire dma_write_addr23_to_bank31      =  (dma__memc__write_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr23_to_bank31       =  (dma__memc__read_address23[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank31   =  dma_write_addr23_to_bank31  & dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank31    =  write_request23_to_bank31   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank31    =  dma_read_addr23_to_bank31   & dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank31     =  read_request23_to_bank31    & memc__dma__read_ready23   ;                                         
  // DMA 24
  wire read_pause24     =  dma__memc__read_pause24   ;  
  // DMA 24, bank0
  wire dma_write_addr24_to_bank0      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr24_to_bank0       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank0   =  dma_write_addr24_to_bank0  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank0    =  write_request24_to_bank0   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank0    =  dma_read_addr24_to_bank0   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank0     =  read_request24_to_bank0    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank1
  wire dma_write_addr24_to_bank1      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr24_to_bank1       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank1   =  dma_write_addr24_to_bank1  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank1    =  write_request24_to_bank1   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank1    =  dma_read_addr24_to_bank1   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank1     =  read_request24_to_bank1    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank2
  wire dma_write_addr24_to_bank2      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr24_to_bank2       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank2   =  dma_write_addr24_to_bank2  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank2    =  write_request24_to_bank2   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank2    =  dma_read_addr24_to_bank2   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank2     =  read_request24_to_bank2    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank3
  wire dma_write_addr24_to_bank3      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr24_to_bank3       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank3   =  dma_write_addr24_to_bank3  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank3    =  write_request24_to_bank3   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank3    =  dma_read_addr24_to_bank3   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank3     =  read_request24_to_bank3    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank4
  wire dma_write_addr24_to_bank4      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr24_to_bank4       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank4   =  dma_write_addr24_to_bank4  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank4    =  write_request24_to_bank4   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank4    =  dma_read_addr24_to_bank4   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank4     =  read_request24_to_bank4    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank5
  wire dma_write_addr24_to_bank5      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr24_to_bank5       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank5   =  dma_write_addr24_to_bank5  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank5    =  write_request24_to_bank5   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank5    =  dma_read_addr24_to_bank5   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank5     =  read_request24_to_bank5    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank6
  wire dma_write_addr24_to_bank6      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr24_to_bank6       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank6   =  dma_write_addr24_to_bank6  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank6    =  write_request24_to_bank6   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank6    =  dma_read_addr24_to_bank6   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank6     =  read_request24_to_bank6    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank7
  wire dma_write_addr24_to_bank7      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr24_to_bank7       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank7   =  dma_write_addr24_to_bank7  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank7    =  write_request24_to_bank7   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank7    =  dma_read_addr24_to_bank7   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank7     =  read_request24_to_bank7    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank8
  wire dma_write_addr24_to_bank8      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr24_to_bank8       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank8   =  dma_write_addr24_to_bank8  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank8    =  write_request24_to_bank8   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank8    =  dma_read_addr24_to_bank8   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank8     =  read_request24_to_bank8    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank9
  wire dma_write_addr24_to_bank9      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr24_to_bank9       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank9   =  dma_write_addr24_to_bank9  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank9    =  write_request24_to_bank9   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank9    =  dma_read_addr24_to_bank9   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank9     =  read_request24_to_bank9    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank10
  wire dma_write_addr24_to_bank10      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr24_to_bank10       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank10   =  dma_write_addr24_to_bank10  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank10    =  write_request24_to_bank10   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank10    =  dma_read_addr24_to_bank10   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank10     =  read_request24_to_bank10    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank11
  wire dma_write_addr24_to_bank11      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr24_to_bank11       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank11   =  dma_write_addr24_to_bank11  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank11    =  write_request24_to_bank11   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank11    =  dma_read_addr24_to_bank11   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank11     =  read_request24_to_bank11    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank12
  wire dma_write_addr24_to_bank12      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr24_to_bank12       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank12   =  dma_write_addr24_to_bank12  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank12    =  write_request24_to_bank12   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank12    =  dma_read_addr24_to_bank12   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank12     =  read_request24_to_bank12    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank13
  wire dma_write_addr24_to_bank13      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr24_to_bank13       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank13   =  dma_write_addr24_to_bank13  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank13    =  write_request24_to_bank13   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank13    =  dma_read_addr24_to_bank13   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank13     =  read_request24_to_bank13    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank14
  wire dma_write_addr24_to_bank14      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr24_to_bank14       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank14   =  dma_write_addr24_to_bank14  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank14    =  write_request24_to_bank14   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank14    =  dma_read_addr24_to_bank14   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank14     =  read_request24_to_bank14    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank15
  wire dma_write_addr24_to_bank15      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr24_to_bank15       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank15   =  dma_write_addr24_to_bank15  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank15    =  write_request24_to_bank15   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank15    =  dma_read_addr24_to_bank15   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank15     =  read_request24_to_bank15    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank16
  wire dma_write_addr24_to_bank16      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr24_to_bank16       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank16   =  dma_write_addr24_to_bank16  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank16    =  write_request24_to_bank16   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank16    =  dma_read_addr24_to_bank16   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank16     =  read_request24_to_bank16    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank17
  wire dma_write_addr24_to_bank17      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr24_to_bank17       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank17   =  dma_write_addr24_to_bank17  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank17    =  write_request24_to_bank17   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank17    =  dma_read_addr24_to_bank17   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank17     =  read_request24_to_bank17    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank18
  wire dma_write_addr24_to_bank18      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr24_to_bank18       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank18   =  dma_write_addr24_to_bank18  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank18    =  write_request24_to_bank18   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank18    =  dma_read_addr24_to_bank18   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank18     =  read_request24_to_bank18    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank19
  wire dma_write_addr24_to_bank19      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr24_to_bank19       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank19   =  dma_write_addr24_to_bank19  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank19    =  write_request24_to_bank19   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank19    =  dma_read_addr24_to_bank19   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank19     =  read_request24_to_bank19    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank20
  wire dma_write_addr24_to_bank20      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr24_to_bank20       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank20   =  dma_write_addr24_to_bank20  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank20    =  write_request24_to_bank20   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank20    =  dma_read_addr24_to_bank20   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank20     =  read_request24_to_bank20    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank21
  wire dma_write_addr24_to_bank21      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr24_to_bank21       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank21   =  dma_write_addr24_to_bank21  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank21    =  write_request24_to_bank21   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank21    =  dma_read_addr24_to_bank21   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank21     =  read_request24_to_bank21    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank22
  wire dma_write_addr24_to_bank22      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr24_to_bank22       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank22   =  dma_write_addr24_to_bank22  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank22    =  write_request24_to_bank22   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank22    =  dma_read_addr24_to_bank22   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank22     =  read_request24_to_bank22    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank23
  wire dma_write_addr24_to_bank23      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr24_to_bank23       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank23   =  dma_write_addr24_to_bank23  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank23    =  write_request24_to_bank23   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank23    =  dma_read_addr24_to_bank23   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank23     =  read_request24_to_bank23    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank24
  wire dma_write_addr24_to_bank24      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr24_to_bank24       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank24   =  dma_write_addr24_to_bank24  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank24    =  write_request24_to_bank24   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank24    =  dma_read_addr24_to_bank24   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank24     =  read_request24_to_bank24    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank25
  wire dma_write_addr24_to_bank25      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr24_to_bank25       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank25   =  dma_write_addr24_to_bank25  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank25    =  write_request24_to_bank25   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank25    =  dma_read_addr24_to_bank25   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank25     =  read_request24_to_bank25    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank26
  wire dma_write_addr24_to_bank26      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr24_to_bank26       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank26   =  dma_write_addr24_to_bank26  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank26    =  write_request24_to_bank26   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank26    =  dma_read_addr24_to_bank26   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank26     =  read_request24_to_bank26    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank27
  wire dma_write_addr24_to_bank27      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr24_to_bank27       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank27   =  dma_write_addr24_to_bank27  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank27    =  write_request24_to_bank27   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank27    =  dma_read_addr24_to_bank27   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank27     =  read_request24_to_bank27    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank28
  wire dma_write_addr24_to_bank28      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr24_to_bank28       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank28   =  dma_write_addr24_to_bank28  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank28    =  write_request24_to_bank28   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank28    =  dma_read_addr24_to_bank28   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank28     =  read_request24_to_bank28    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank29
  wire dma_write_addr24_to_bank29      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr24_to_bank29       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank29   =  dma_write_addr24_to_bank29  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank29    =  write_request24_to_bank29   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank29    =  dma_read_addr24_to_bank29   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank29     =  read_request24_to_bank29    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank30
  wire dma_write_addr24_to_bank30      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr24_to_bank30       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank30   =  dma_write_addr24_to_bank30  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank30    =  write_request24_to_bank30   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank30    =  dma_read_addr24_to_bank30   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank30     =  read_request24_to_bank30    & memc__dma__read_ready24   ;                                         
  // DMA 24, bank31
  wire dma_write_addr24_to_bank31      =  (dma__memc__write_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr24_to_bank31       =  (dma__memc__read_address24[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank31   =  dma_write_addr24_to_bank31  & dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank31    =  write_request24_to_bank31   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank31    =  dma_read_addr24_to_bank31   & dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank31     =  read_request24_to_bank31    & memc__dma__read_ready24   ;                                         
  // DMA 25
  wire read_pause25     =  dma__memc__read_pause25   ;  
  // DMA 25, bank0
  wire dma_write_addr25_to_bank0      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr25_to_bank0       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank0   =  dma_write_addr25_to_bank0  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank0    =  write_request25_to_bank0   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank0    =  dma_read_addr25_to_bank0   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank0     =  read_request25_to_bank0    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank1
  wire dma_write_addr25_to_bank1      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr25_to_bank1       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank1   =  dma_write_addr25_to_bank1  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank1    =  write_request25_to_bank1   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank1    =  dma_read_addr25_to_bank1   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank1     =  read_request25_to_bank1    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank2
  wire dma_write_addr25_to_bank2      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr25_to_bank2       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank2   =  dma_write_addr25_to_bank2  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank2    =  write_request25_to_bank2   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank2    =  dma_read_addr25_to_bank2   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank2     =  read_request25_to_bank2    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank3
  wire dma_write_addr25_to_bank3      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr25_to_bank3       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank3   =  dma_write_addr25_to_bank3  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank3    =  write_request25_to_bank3   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank3    =  dma_read_addr25_to_bank3   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank3     =  read_request25_to_bank3    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank4
  wire dma_write_addr25_to_bank4      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr25_to_bank4       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank4   =  dma_write_addr25_to_bank4  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank4    =  write_request25_to_bank4   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank4    =  dma_read_addr25_to_bank4   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank4     =  read_request25_to_bank4    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank5
  wire dma_write_addr25_to_bank5      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr25_to_bank5       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank5   =  dma_write_addr25_to_bank5  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank5    =  write_request25_to_bank5   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank5    =  dma_read_addr25_to_bank5   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank5     =  read_request25_to_bank5    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank6
  wire dma_write_addr25_to_bank6      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr25_to_bank6       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank6   =  dma_write_addr25_to_bank6  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank6    =  write_request25_to_bank6   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank6    =  dma_read_addr25_to_bank6   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank6     =  read_request25_to_bank6    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank7
  wire dma_write_addr25_to_bank7      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr25_to_bank7       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank7   =  dma_write_addr25_to_bank7  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank7    =  write_request25_to_bank7   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank7    =  dma_read_addr25_to_bank7   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank7     =  read_request25_to_bank7    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank8
  wire dma_write_addr25_to_bank8      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr25_to_bank8       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank8   =  dma_write_addr25_to_bank8  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank8    =  write_request25_to_bank8   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank8    =  dma_read_addr25_to_bank8   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank8     =  read_request25_to_bank8    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank9
  wire dma_write_addr25_to_bank9      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr25_to_bank9       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank9   =  dma_write_addr25_to_bank9  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank9    =  write_request25_to_bank9   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank9    =  dma_read_addr25_to_bank9   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank9     =  read_request25_to_bank9    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank10
  wire dma_write_addr25_to_bank10      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr25_to_bank10       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank10   =  dma_write_addr25_to_bank10  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank10    =  write_request25_to_bank10   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank10    =  dma_read_addr25_to_bank10   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank10     =  read_request25_to_bank10    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank11
  wire dma_write_addr25_to_bank11      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr25_to_bank11       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank11   =  dma_write_addr25_to_bank11  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank11    =  write_request25_to_bank11   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank11    =  dma_read_addr25_to_bank11   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank11     =  read_request25_to_bank11    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank12
  wire dma_write_addr25_to_bank12      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr25_to_bank12       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank12   =  dma_write_addr25_to_bank12  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank12    =  write_request25_to_bank12   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank12    =  dma_read_addr25_to_bank12   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank12     =  read_request25_to_bank12    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank13
  wire dma_write_addr25_to_bank13      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr25_to_bank13       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank13   =  dma_write_addr25_to_bank13  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank13    =  write_request25_to_bank13   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank13    =  dma_read_addr25_to_bank13   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank13     =  read_request25_to_bank13    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank14
  wire dma_write_addr25_to_bank14      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr25_to_bank14       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank14   =  dma_write_addr25_to_bank14  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank14    =  write_request25_to_bank14   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank14    =  dma_read_addr25_to_bank14   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank14     =  read_request25_to_bank14    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank15
  wire dma_write_addr25_to_bank15      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr25_to_bank15       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank15   =  dma_write_addr25_to_bank15  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank15    =  write_request25_to_bank15   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank15    =  dma_read_addr25_to_bank15   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank15     =  read_request25_to_bank15    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank16
  wire dma_write_addr25_to_bank16      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr25_to_bank16       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank16   =  dma_write_addr25_to_bank16  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank16    =  write_request25_to_bank16   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank16    =  dma_read_addr25_to_bank16   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank16     =  read_request25_to_bank16    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank17
  wire dma_write_addr25_to_bank17      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr25_to_bank17       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank17   =  dma_write_addr25_to_bank17  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank17    =  write_request25_to_bank17   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank17    =  dma_read_addr25_to_bank17   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank17     =  read_request25_to_bank17    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank18
  wire dma_write_addr25_to_bank18      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr25_to_bank18       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank18   =  dma_write_addr25_to_bank18  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank18    =  write_request25_to_bank18   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank18    =  dma_read_addr25_to_bank18   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank18     =  read_request25_to_bank18    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank19
  wire dma_write_addr25_to_bank19      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr25_to_bank19       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank19   =  dma_write_addr25_to_bank19  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank19    =  write_request25_to_bank19   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank19    =  dma_read_addr25_to_bank19   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank19     =  read_request25_to_bank19    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank20
  wire dma_write_addr25_to_bank20      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr25_to_bank20       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank20   =  dma_write_addr25_to_bank20  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank20    =  write_request25_to_bank20   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank20    =  dma_read_addr25_to_bank20   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank20     =  read_request25_to_bank20    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank21
  wire dma_write_addr25_to_bank21      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr25_to_bank21       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank21   =  dma_write_addr25_to_bank21  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank21    =  write_request25_to_bank21   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank21    =  dma_read_addr25_to_bank21   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank21     =  read_request25_to_bank21    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank22
  wire dma_write_addr25_to_bank22      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr25_to_bank22       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank22   =  dma_write_addr25_to_bank22  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank22    =  write_request25_to_bank22   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank22    =  dma_read_addr25_to_bank22   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank22     =  read_request25_to_bank22    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank23
  wire dma_write_addr25_to_bank23      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr25_to_bank23       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank23   =  dma_write_addr25_to_bank23  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank23    =  write_request25_to_bank23   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank23    =  dma_read_addr25_to_bank23   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank23     =  read_request25_to_bank23    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank24
  wire dma_write_addr25_to_bank24      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr25_to_bank24       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank24   =  dma_write_addr25_to_bank24  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank24    =  write_request25_to_bank24   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank24    =  dma_read_addr25_to_bank24   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank24     =  read_request25_to_bank24    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank25
  wire dma_write_addr25_to_bank25      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr25_to_bank25       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank25   =  dma_write_addr25_to_bank25  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank25    =  write_request25_to_bank25   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank25    =  dma_read_addr25_to_bank25   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank25     =  read_request25_to_bank25    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank26
  wire dma_write_addr25_to_bank26      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr25_to_bank26       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank26   =  dma_write_addr25_to_bank26  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank26    =  write_request25_to_bank26   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank26    =  dma_read_addr25_to_bank26   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank26     =  read_request25_to_bank26    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank27
  wire dma_write_addr25_to_bank27      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr25_to_bank27       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank27   =  dma_write_addr25_to_bank27  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank27    =  write_request25_to_bank27   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank27    =  dma_read_addr25_to_bank27   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank27     =  read_request25_to_bank27    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank28
  wire dma_write_addr25_to_bank28      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr25_to_bank28       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank28   =  dma_write_addr25_to_bank28  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank28    =  write_request25_to_bank28   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank28    =  dma_read_addr25_to_bank28   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank28     =  read_request25_to_bank28    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank29
  wire dma_write_addr25_to_bank29      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr25_to_bank29       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank29   =  dma_write_addr25_to_bank29  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank29    =  write_request25_to_bank29   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank29    =  dma_read_addr25_to_bank29   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank29     =  read_request25_to_bank29    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank30
  wire dma_write_addr25_to_bank30      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr25_to_bank30       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank30   =  dma_write_addr25_to_bank30  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank30    =  write_request25_to_bank30   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank30    =  dma_read_addr25_to_bank30   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank30     =  read_request25_to_bank30    & memc__dma__read_ready25   ;                                         
  // DMA 25, bank31
  wire dma_write_addr25_to_bank31      =  (dma__memc__write_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr25_to_bank31       =  (dma__memc__read_address25[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank31   =  dma_write_addr25_to_bank31  & dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank31    =  write_request25_to_bank31   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank31    =  dma_read_addr25_to_bank31   & dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank31     =  read_request25_to_bank31    & memc__dma__read_ready25   ;                                         
  // DMA 26
  wire read_pause26     =  dma__memc__read_pause26   ;  
  // DMA 26, bank0
  wire dma_write_addr26_to_bank0      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr26_to_bank0       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank0   =  dma_write_addr26_to_bank0  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank0    =  write_request26_to_bank0   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank0    =  dma_read_addr26_to_bank0   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank0     =  read_request26_to_bank0    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank1
  wire dma_write_addr26_to_bank1      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr26_to_bank1       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank1   =  dma_write_addr26_to_bank1  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank1    =  write_request26_to_bank1   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank1    =  dma_read_addr26_to_bank1   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank1     =  read_request26_to_bank1    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank2
  wire dma_write_addr26_to_bank2      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr26_to_bank2       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank2   =  dma_write_addr26_to_bank2  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank2    =  write_request26_to_bank2   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank2    =  dma_read_addr26_to_bank2   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank2     =  read_request26_to_bank2    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank3
  wire dma_write_addr26_to_bank3      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr26_to_bank3       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank3   =  dma_write_addr26_to_bank3  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank3    =  write_request26_to_bank3   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank3    =  dma_read_addr26_to_bank3   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank3     =  read_request26_to_bank3    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank4
  wire dma_write_addr26_to_bank4      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr26_to_bank4       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank4   =  dma_write_addr26_to_bank4  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank4    =  write_request26_to_bank4   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank4    =  dma_read_addr26_to_bank4   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank4     =  read_request26_to_bank4    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank5
  wire dma_write_addr26_to_bank5      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr26_to_bank5       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank5   =  dma_write_addr26_to_bank5  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank5    =  write_request26_to_bank5   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank5    =  dma_read_addr26_to_bank5   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank5     =  read_request26_to_bank5    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank6
  wire dma_write_addr26_to_bank6      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr26_to_bank6       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank6   =  dma_write_addr26_to_bank6  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank6    =  write_request26_to_bank6   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank6    =  dma_read_addr26_to_bank6   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank6     =  read_request26_to_bank6    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank7
  wire dma_write_addr26_to_bank7      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr26_to_bank7       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank7   =  dma_write_addr26_to_bank7  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank7    =  write_request26_to_bank7   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank7    =  dma_read_addr26_to_bank7   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank7     =  read_request26_to_bank7    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank8
  wire dma_write_addr26_to_bank8      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr26_to_bank8       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank8   =  dma_write_addr26_to_bank8  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank8    =  write_request26_to_bank8   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank8    =  dma_read_addr26_to_bank8   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank8     =  read_request26_to_bank8    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank9
  wire dma_write_addr26_to_bank9      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr26_to_bank9       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank9   =  dma_write_addr26_to_bank9  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank9    =  write_request26_to_bank9   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank9    =  dma_read_addr26_to_bank9   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank9     =  read_request26_to_bank9    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank10
  wire dma_write_addr26_to_bank10      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr26_to_bank10       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank10   =  dma_write_addr26_to_bank10  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank10    =  write_request26_to_bank10   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank10    =  dma_read_addr26_to_bank10   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank10     =  read_request26_to_bank10    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank11
  wire dma_write_addr26_to_bank11      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr26_to_bank11       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank11   =  dma_write_addr26_to_bank11  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank11    =  write_request26_to_bank11   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank11    =  dma_read_addr26_to_bank11   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank11     =  read_request26_to_bank11    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank12
  wire dma_write_addr26_to_bank12      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr26_to_bank12       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank12   =  dma_write_addr26_to_bank12  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank12    =  write_request26_to_bank12   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank12    =  dma_read_addr26_to_bank12   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank12     =  read_request26_to_bank12    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank13
  wire dma_write_addr26_to_bank13      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr26_to_bank13       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank13   =  dma_write_addr26_to_bank13  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank13    =  write_request26_to_bank13   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank13    =  dma_read_addr26_to_bank13   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank13     =  read_request26_to_bank13    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank14
  wire dma_write_addr26_to_bank14      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr26_to_bank14       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank14   =  dma_write_addr26_to_bank14  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank14    =  write_request26_to_bank14   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank14    =  dma_read_addr26_to_bank14   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank14     =  read_request26_to_bank14    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank15
  wire dma_write_addr26_to_bank15      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr26_to_bank15       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank15   =  dma_write_addr26_to_bank15  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank15    =  write_request26_to_bank15   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank15    =  dma_read_addr26_to_bank15   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank15     =  read_request26_to_bank15    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank16
  wire dma_write_addr26_to_bank16      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr26_to_bank16       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank16   =  dma_write_addr26_to_bank16  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank16    =  write_request26_to_bank16   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank16    =  dma_read_addr26_to_bank16   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank16     =  read_request26_to_bank16    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank17
  wire dma_write_addr26_to_bank17      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr26_to_bank17       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank17   =  dma_write_addr26_to_bank17  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank17    =  write_request26_to_bank17   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank17    =  dma_read_addr26_to_bank17   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank17     =  read_request26_to_bank17    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank18
  wire dma_write_addr26_to_bank18      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr26_to_bank18       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank18   =  dma_write_addr26_to_bank18  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank18    =  write_request26_to_bank18   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank18    =  dma_read_addr26_to_bank18   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank18     =  read_request26_to_bank18    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank19
  wire dma_write_addr26_to_bank19      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr26_to_bank19       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank19   =  dma_write_addr26_to_bank19  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank19    =  write_request26_to_bank19   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank19    =  dma_read_addr26_to_bank19   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank19     =  read_request26_to_bank19    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank20
  wire dma_write_addr26_to_bank20      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr26_to_bank20       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank20   =  dma_write_addr26_to_bank20  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank20    =  write_request26_to_bank20   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank20    =  dma_read_addr26_to_bank20   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank20     =  read_request26_to_bank20    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank21
  wire dma_write_addr26_to_bank21      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr26_to_bank21       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank21   =  dma_write_addr26_to_bank21  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank21    =  write_request26_to_bank21   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank21    =  dma_read_addr26_to_bank21   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank21     =  read_request26_to_bank21    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank22
  wire dma_write_addr26_to_bank22      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr26_to_bank22       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank22   =  dma_write_addr26_to_bank22  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank22    =  write_request26_to_bank22   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank22    =  dma_read_addr26_to_bank22   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank22     =  read_request26_to_bank22    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank23
  wire dma_write_addr26_to_bank23      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr26_to_bank23       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank23   =  dma_write_addr26_to_bank23  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank23    =  write_request26_to_bank23   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank23    =  dma_read_addr26_to_bank23   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank23     =  read_request26_to_bank23    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank24
  wire dma_write_addr26_to_bank24      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr26_to_bank24       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank24   =  dma_write_addr26_to_bank24  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank24    =  write_request26_to_bank24   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank24    =  dma_read_addr26_to_bank24   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank24     =  read_request26_to_bank24    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank25
  wire dma_write_addr26_to_bank25      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr26_to_bank25       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank25   =  dma_write_addr26_to_bank25  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank25    =  write_request26_to_bank25   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank25    =  dma_read_addr26_to_bank25   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank25     =  read_request26_to_bank25    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank26
  wire dma_write_addr26_to_bank26      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr26_to_bank26       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank26   =  dma_write_addr26_to_bank26  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank26    =  write_request26_to_bank26   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank26    =  dma_read_addr26_to_bank26   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank26     =  read_request26_to_bank26    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank27
  wire dma_write_addr26_to_bank27      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr26_to_bank27       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank27   =  dma_write_addr26_to_bank27  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank27    =  write_request26_to_bank27   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank27    =  dma_read_addr26_to_bank27   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank27     =  read_request26_to_bank27    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank28
  wire dma_write_addr26_to_bank28      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr26_to_bank28       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank28   =  dma_write_addr26_to_bank28  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank28    =  write_request26_to_bank28   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank28    =  dma_read_addr26_to_bank28   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank28     =  read_request26_to_bank28    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank29
  wire dma_write_addr26_to_bank29      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr26_to_bank29       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank29   =  dma_write_addr26_to_bank29  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank29    =  write_request26_to_bank29   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank29    =  dma_read_addr26_to_bank29   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank29     =  read_request26_to_bank29    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank30
  wire dma_write_addr26_to_bank30      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr26_to_bank30       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank30   =  dma_write_addr26_to_bank30  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank30    =  write_request26_to_bank30   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank30    =  dma_read_addr26_to_bank30   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank30     =  read_request26_to_bank30    & memc__dma__read_ready26   ;                                         
  // DMA 26, bank31
  wire dma_write_addr26_to_bank31      =  (dma__memc__write_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr26_to_bank31       =  (dma__memc__read_address26[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank31   =  dma_write_addr26_to_bank31  & dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank31    =  write_request26_to_bank31   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank31    =  dma_read_addr26_to_bank31   & dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank31     =  read_request26_to_bank31    & memc__dma__read_ready26   ;                                         
  // DMA 27
  wire read_pause27     =  dma__memc__read_pause27   ;  
  // DMA 27, bank0
  wire dma_write_addr27_to_bank0      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr27_to_bank0       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank0   =  dma_write_addr27_to_bank0  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank0    =  write_request27_to_bank0   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank0    =  dma_read_addr27_to_bank0   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank0     =  read_request27_to_bank0    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank1
  wire dma_write_addr27_to_bank1      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr27_to_bank1       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank1   =  dma_write_addr27_to_bank1  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank1    =  write_request27_to_bank1   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank1    =  dma_read_addr27_to_bank1   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank1     =  read_request27_to_bank1    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank2
  wire dma_write_addr27_to_bank2      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr27_to_bank2       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank2   =  dma_write_addr27_to_bank2  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank2    =  write_request27_to_bank2   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank2    =  dma_read_addr27_to_bank2   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank2     =  read_request27_to_bank2    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank3
  wire dma_write_addr27_to_bank3      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr27_to_bank3       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank3   =  dma_write_addr27_to_bank3  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank3    =  write_request27_to_bank3   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank3    =  dma_read_addr27_to_bank3   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank3     =  read_request27_to_bank3    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank4
  wire dma_write_addr27_to_bank4      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr27_to_bank4       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank4   =  dma_write_addr27_to_bank4  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank4    =  write_request27_to_bank4   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank4    =  dma_read_addr27_to_bank4   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank4     =  read_request27_to_bank4    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank5
  wire dma_write_addr27_to_bank5      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr27_to_bank5       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank5   =  dma_write_addr27_to_bank5  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank5    =  write_request27_to_bank5   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank5    =  dma_read_addr27_to_bank5   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank5     =  read_request27_to_bank5    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank6
  wire dma_write_addr27_to_bank6      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr27_to_bank6       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank6   =  dma_write_addr27_to_bank6  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank6    =  write_request27_to_bank6   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank6    =  dma_read_addr27_to_bank6   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank6     =  read_request27_to_bank6    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank7
  wire dma_write_addr27_to_bank7      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr27_to_bank7       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank7   =  dma_write_addr27_to_bank7  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank7    =  write_request27_to_bank7   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank7    =  dma_read_addr27_to_bank7   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank7     =  read_request27_to_bank7    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank8
  wire dma_write_addr27_to_bank8      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr27_to_bank8       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank8   =  dma_write_addr27_to_bank8  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank8    =  write_request27_to_bank8   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank8    =  dma_read_addr27_to_bank8   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank8     =  read_request27_to_bank8    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank9
  wire dma_write_addr27_to_bank9      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr27_to_bank9       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank9   =  dma_write_addr27_to_bank9  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank9    =  write_request27_to_bank9   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank9    =  dma_read_addr27_to_bank9   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank9     =  read_request27_to_bank9    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank10
  wire dma_write_addr27_to_bank10      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr27_to_bank10       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank10   =  dma_write_addr27_to_bank10  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank10    =  write_request27_to_bank10   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank10    =  dma_read_addr27_to_bank10   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank10     =  read_request27_to_bank10    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank11
  wire dma_write_addr27_to_bank11      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr27_to_bank11       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank11   =  dma_write_addr27_to_bank11  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank11    =  write_request27_to_bank11   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank11    =  dma_read_addr27_to_bank11   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank11     =  read_request27_to_bank11    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank12
  wire dma_write_addr27_to_bank12      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr27_to_bank12       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank12   =  dma_write_addr27_to_bank12  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank12    =  write_request27_to_bank12   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank12    =  dma_read_addr27_to_bank12   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank12     =  read_request27_to_bank12    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank13
  wire dma_write_addr27_to_bank13      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr27_to_bank13       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank13   =  dma_write_addr27_to_bank13  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank13    =  write_request27_to_bank13   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank13    =  dma_read_addr27_to_bank13   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank13     =  read_request27_to_bank13    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank14
  wire dma_write_addr27_to_bank14      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr27_to_bank14       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank14   =  dma_write_addr27_to_bank14  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank14    =  write_request27_to_bank14   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank14    =  dma_read_addr27_to_bank14   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank14     =  read_request27_to_bank14    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank15
  wire dma_write_addr27_to_bank15      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr27_to_bank15       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank15   =  dma_write_addr27_to_bank15  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank15    =  write_request27_to_bank15   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank15    =  dma_read_addr27_to_bank15   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank15     =  read_request27_to_bank15    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank16
  wire dma_write_addr27_to_bank16      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr27_to_bank16       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank16   =  dma_write_addr27_to_bank16  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank16    =  write_request27_to_bank16   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank16    =  dma_read_addr27_to_bank16   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank16     =  read_request27_to_bank16    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank17
  wire dma_write_addr27_to_bank17      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr27_to_bank17       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank17   =  dma_write_addr27_to_bank17  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank17    =  write_request27_to_bank17   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank17    =  dma_read_addr27_to_bank17   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank17     =  read_request27_to_bank17    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank18
  wire dma_write_addr27_to_bank18      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr27_to_bank18       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank18   =  dma_write_addr27_to_bank18  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank18    =  write_request27_to_bank18   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank18    =  dma_read_addr27_to_bank18   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank18     =  read_request27_to_bank18    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank19
  wire dma_write_addr27_to_bank19      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr27_to_bank19       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank19   =  dma_write_addr27_to_bank19  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank19    =  write_request27_to_bank19   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank19    =  dma_read_addr27_to_bank19   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank19     =  read_request27_to_bank19    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank20
  wire dma_write_addr27_to_bank20      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr27_to_bank20       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank20   =  dma_write_addr27_to_bank20  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank20    =  write_request27_to_bank20   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank20    =  dma_read_addr27_to_bank20   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank20     =  read_request27_to_bank20    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank21
  wire dma_write_addr27_to_bank21      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr27_to_bank21       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank21   =  dma_write_addr27_to_bank21  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank21    =  write_request27_to_bank21   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank21    =  dma_read_addr27_to_bank21   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank21     =  read_request27_to_bank21    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank22
  wire dma_write_addr27_to_bank22      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr27_to_bank22       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank22   =  dma_write_addr27_to_bank22  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank22    =  write_request27_to_bank22   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank22    =  dma_read_addr27_to_bank22   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank22     =  read_request27_to_bank22    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank23
  wire dma_write_addr27_to_bank23      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr27_to_bank23       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank23   =  dma_write_addr27_to_bank23  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank23    =  write_request27_to_bank23   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank23    =  dma_read_addr27_to_bank23   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank23     =  read_request27_to_bank23    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank24
  wire dma_write_addr27_to_bank24      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr27_to_bank24       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank24   =  dma_write_addr27_to_bank24  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank24    =  write_request27_to_bank24   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank24    =  dma_read_addr27_to_bank24   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank24     =  read_request27_to_bank24    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank25
  wire dma_write_addr27_to_bank25      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr27_to_bank25       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank25   =  dma_write_addr27_to_bank25  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank25    =  write_request27_to_bank25   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank25    =  dma_read_addr27_to_bank25   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank25     =  read_request27_to_bank25    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank26
  wire dma_write_addr27_to_bank26      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr27_to_bank26       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank26   =  dma_write_addr27_to_bank26  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank26    =  write_request27_to_bank26   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank26    =  dma_read_addr27_to_bank26   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank26     =  read_request27_to_bank26    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank27
  wire dma_write_addr27_to_bank27      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr27_to_bank27       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank27   =  dma_write_addr27_to_bank27  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank27    =  write_request27_to_bank27   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank27    =  dma_read_addr27_to_bank27   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank27     =  read_request27_to_bank27    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank28
  wire dma_write_addr27_to_bank28      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr27_to_bank28       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank28   =  dma_write_addr27_to_bank28  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank28    =  write_request27_to_bank28   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank28    =  dma_read_addr27_to_bank28   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank28     =  read_request27_to_bank28    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank29
  wire dma_write_addr27_to_bank29      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr27_to_bank29       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank29   =  dma_write_addr27_to_bank29  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank29    =  write_request27_to_bank29   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank29    =  dma_read_addr27_to_bank29   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank29     =  read_request27_to_bank29    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank30
  wire dma_write_addr27_to_bank30      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr27_to_bank30       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank30   =  dma_write_addr27_to_bank30  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank30    =  write_request27_to_bank30   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank30    =  dma_read_addr27_to_bank30   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank30     =  read_request27_to_bank30    & memc__dma__read_ready27   ;                                         
  // DMA 27, bank31
  wire dma_write_addr27_to_bank31      =  (dma__memc__write_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr27_to_bank31       =  (dma__memc__read_address27[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank31   =  dma_write_addr27_to_bank31  & dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank31    =  write_request27_to_bank31   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank31    =  dma_read_addr27_to_bank31   & dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank31     =  read_request27_to_bank31    & memc__dma__read_ready27   ;                                         
  // DMA 28
  wire read_pause28     =  dma__memc__read_pause28   ;  
  // DMA 28, bank0
  wire dma_write_addr28_to_bank0      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr28_to_bank0       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank0   =  dma_write_addr28_to_bank0  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank0    =  write_request28_to_bank0   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank0    =  dma_read_addr28_to_bank0   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank0     =  read_request28_to_bank0    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank1
  wire dma_write_addr28_to_bank1      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr28_to_bank1       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank1   =  dma_write_addr28_to_bank1  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank1    =  write_request28_to_bank1   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank1    =  dma_read_addr28_to_bank1   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank1     =  read_request28_to_bank1    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank2
  wire dma_write_addr28_to_bank2      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr28_to_bank2       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank2   =  dma_write_addr28_to_bank2  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank2    =  write_request28_to_bank2   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank2    =  dma_read_addr28_to_bank2   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank2     =  read_request28_to_bank2    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank3
  wire dma_write_addr28_to_bank3      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr28_to_bank3       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank3   =  dma_write_addr28_to_bank3  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank3    =  write_request28_to_bank3   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank3    =  dma_read_addr28_to_bank3   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank3     =  read_request28_to_bank3    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank4
  wire dma_write_addr28_to_bank4      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr28_to_bank4       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank4   =  dma_write_addr28_to_bank4  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank4    =  write_request28_to_bank4   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank4    =  dma_read_addr28_to_bank4   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank4     =  read_request28_to_bank4    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank5
  wire dma_write_addr28_to_bank5      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr28_to_bank5       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank5   =  dma_write_addr28_to_bank5  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank5    =  write_request28_to_bank5   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank5    =  dma_read_addr28_to_bank5   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank5     =  read_request28_to_bank5    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank6
  wire dma_write_addr28_to_bank6      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr28_to_bank6       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank6   =  dma_write_addr28_to_bank6  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank6    =  write_request28_to_bank6   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank6    =  dma_read_addr28_to_bank6   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank6     =  read_request28_to_bank6    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank7
  wire dma_write_addr28_to_bank7      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr28_to_bank7       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank7   =  dma_write_addr28_to_bank7  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank7    =  write_request28_to_bank7   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank7    =  dma_read_addr28_to_bank7   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank7     =  read_request28_to_bank7    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank8
  wire dma_write_addr28_to_bank8      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr28_to_bank8       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank8   =  dma_write_addr28_to_bank8  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank8    =  write_request28_to_bank8   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank8    =  dma_read_addr28_to_bank8   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank8     =  read_request28_to_bank8    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank9
  wire dma_write_addr28_to_bank9      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr28_to_bank9       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank9   =  dma_write_addr28_to_bank9  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank9    =  write_request28_to_bank9   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank9    =  dma_read_addr28_to_bank9   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank9     =  read_request28_to_bank9    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank10
  wire dma_write_addr28_to_bank10      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr28_to_bank10       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank10   =  dma_write_addr28_to_bank10  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank10    =  write_request28_to_bank10   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank10    =  dma_read_addr28_to_bank10   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank10     =  read_request28_to_bank10    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank11
  wire dma_write_addr28_to_bank11      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr28_to_bank11       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank11   =  dma_write_addr28_to_bank11  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank11    =  write_request28_to_bank11   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank11    =  dma_read_addr28_to_bank11   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank11     =  read_request28_to_bank11    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank12
  wire dma_write_addr28_to_bank12      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr28_to_bank12       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank12   =  dma_write_addr28_to_bank12  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank12    =  write_request28_to_bank12   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank12    =  dma_read_addr28_to_bank12   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank12     =  read_request28_to_bank12    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank13
  wire dma_write_addr28_to_bank13      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr28_to_bank13       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank13   =  dma_write_addr28_to_bank13  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank13    =  write_request28_to_bank13   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank13    =  dma_read_addr28_to_bank13   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank13     =  read_request28_to_bank13    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank14
  wire dma_write_addr28_to_bank14      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr28_to_bank14       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank14   =  dma_write_addr28_to_bank14  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank14    =  write_request28_to_bank14   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank14    =  dma_read_addr28_to_bank14   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank14     =  read_request28_to_bank14    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank15
  wire dma_write_addr28_to_bank15      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr28_to_bank15       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank15   =  dma_write_addr28_to_bank15  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank15    =  write_request28_to_bank15   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank15    =  dma_read_addr28_to_bank15   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank15     =  read_request28_to_bank15    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank16
  wire dma_write_addr28_to_bank16      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr28_to_bank16       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank16   =  dma_write_addr28_to_bank16  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank16    =  write_request28_to_bank16   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank16    =  dma_read_addr28_to_bank16   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank16     =  read_request28_to_bank16    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank17
  wire dma_write_addr28_to_bank17      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr28_to_bank17       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank17   =  dma_write_addr28_to_bank17  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank17    =  write_request28_to_bank17   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank17    =  dma_read_addr28_to_bank17   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank17     =  read_request28_to_bank17    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank18
  wire dma_write_addr28_to_bank18      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr28_to_bank18       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank18   =  dma_write_addr28_to_bank18  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank18    =  write_request28_to_bank18   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank18    =  dma_read_addr28_to_bank18   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank18     =  read_request28_to_bank18    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank19
  wire dma_write_addr28_to_bank19      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr28_to_bank19       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank19   =  dma_write_addr28_to_bank19  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank19    =  write_request28_to_bank19   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank19    =  dma_read_addr28_to_bank19   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank19     =  read_request28_to_bank19    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank20
  wire dma_write_addr28_to_bank20      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr28_to_bank20       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank20   =  dma_write_addr28_to_bank20  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank20    =  write_request28_to_bank20   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank20    =  dma_read_addr28_to_bank20   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank20     =  read_request28_to_bank20    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank21
  wire dma_write_addr28_to_bank21      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr28_to_bank21       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank21   =  dma_write_addr28_to_bank21  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank21    =  write_request28_to_bank21   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank21    =  dma_read_addr28_to_bank21   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank21     =  read_request28_to_bank21    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank22
  wire dma_write_addr28_to_bank22      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr28_to_bank22       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank22   =  dma_write_addr28_to_bank22  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank22    =  write_request28_to_bank22   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank22    =  dma_read_addr28_to_bank22   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank22     =  read_request28_to_bank22    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank23
  wire dma_write_addr28_to_bank23      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr28_to_bank23       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank23   =  dma_write_addr28_to_bank23  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank23    =  write_request28_to_bank23   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank23    =  dma_read_addr28_to_bank23   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank23     =  read_request28_to_bank23    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank24
  wire dma_write_addr28_to_bank24      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr28_to_bank24       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank24   =  dma_write_addr28_to_bank24  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank24    =  write_request28_to_bank24   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank24    =  dma_read_addr28_to_bank24   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank24     =  read_request28_to_bank24    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank25
  wire dma_write_addr28_to_bank25      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr28_to_bank25       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank25   =  dma_write_addr28_to_bank25  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank25    =  write_request28_to_bank25   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank25    =  dma_read_addr28_to_bank25   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank25     =  read_request28_to_bank25    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank26
  wire dma_write_addr28_to_bank26      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr28_to_bank26       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank26   =  dma_write_addr28_to_bank26  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank26    =  write_request28_to_bank26   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank26    =  dma_read_addr28_to_bank26   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank26     =  read_request28_to_bank26    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank27
  wire dma_write_addr28_to_bank27      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr28_to_bank27       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank27   =  dma_write_addr28_to_bank27  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank27    =  write_request28_to_bank27   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank27    =  dma_read_addr28_to_bank27   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank27     =  read_request28_to_bank27    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank28
  wire dma_write_addr28_to_bank28      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr28_to_bank28       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank28   =  dma_write_addr28_to_bank28  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank28    =  write_request28_to_bank28   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank28    =  dma_read_addr28_to_bank28   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank28     =  read_request28_to_bank28    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank29
  wire dma_write_addr28_to_bank29      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr28_to_bank29       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank29   =  dma_write_addr28_to_bank29  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank29    =  write_request28_to_bank29   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank29    =  dma_read_addr28_to_bank29   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank29     =  read_request28_to_bank29    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank30
  wire dma_write_addr28_to_bank30      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr28_to_bank30       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank30   =  dma_write_addr28_to_bank30  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank30    =  write_request28_to_bank30   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank30    =  dma_read_addr28_to_bank30   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank30     =  read_request28_to_bank30    & memc__dma__read_ready28   ;                                         
  // DMA 28, bank31
  wire dma_write_addr28_to_bank31      =  (dma__memc__write_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr28_to_bank31       =  (dma__memc__read_address28[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank31   =  dma_write_addr28_to_bank31  & dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank31    =  write_request28_to_bank31   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank31    =  dma_read_addr28_to_bank31   & dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank31     =  read_request28_to_bank31    & memc__dma__read_ready28   ;                                         
  // DMA 29
  wire read_pause29     =  dma__memc__read_pause29   ;  
  // DMA 29, bank0
  wire dma_write_addr29_to_bank0      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr29_to_bank0       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank0   =  dma_write_addr29_to_bank0  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank0    =  write_request29_to_bank0   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank0    =  dma_read_addr29_to_bank0   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank0     =  read_request29_to_bank0    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank1
  wire dma_write_addr29_to_bank1      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr29_to_bank1       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank1   =  dma_write_addr29_to_bank1  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank1    =  write_request29_to_bank1   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank1    =  dma_read_addr29_to_bank1   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank1     =  read_request29_to_bank1    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank2
  wire dma_write_addr29_to_bank2      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr29_to_bank2       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank2   =  dma_write_addr29_to_bank2  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank2    =  write_request29_to_bank2   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank2    =  dma_read_addr29_to_bank2   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank2     =  read_request29_to_bank2    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank3
  wire dma_write_addr29_to_bank3      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr29_to_bank3       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank3   =  dma_write_addr29_to_bank3  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank3    =  write_request29_to_bank3   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank3    =  dma_read_addr29_to_bank3   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank3     =  read_request29_to_bank3    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank4
  wire dma_write_addr29_to_bank4      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr29_to_bank4       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank4   =  dma_write_addr29_to_bank4  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank4    =  write_request29_to_bank4   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank4    =  dma_read_addr29_to_bank4   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank4     =  read_request29_to_bank4    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank5
  wire dma_write_addr29_to_bank5      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr29_to_bank5       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank5   =  dma_write_addr29_to_bank5  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank5    =  write_request29_to_bank5   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank5    =  dma_read_addr29_to_bank5   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank5     =  read_request29_to_bank5    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank6
  wire dma_write_addr29_to_bank6      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr29_to_bank6       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank6   =  dma_write_addr29_to_bank6  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank6    =  write_request29_to_bank6   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank6    =  dma_read_addr29_to_bank6   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank6     =  read_request29_to_bank6    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank7
  wire dma_write_addr29_to_bank7      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr29_to_bank7       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank7   =  dma_write_addr29_to_bank7  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank7    =  write_request29_to_bank7   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank7    =  dma_read_addr29_to_bank7   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank7     =  read_request29_to_bank7    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank8
  wire dma_write_addr29_to_bank8      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr29_to_bank8       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank8   =  dma_write_addr29_to_bank8  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank8    =  write_request29_to_bank8   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank8    =  dma_read_addr29_to_bank8   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank8     =  read_request29_to_bank8    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank9
  wire dma_write_addr29_to_bank9      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr29_to_bank9       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank9   =  dma_write_addr29_to_bank9  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank9    =  write_request29_to_bank9   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank9    =  dma_read_addr29_to_bank9   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank9     =  read_request29_to_bank9    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank10
  wire dma_write_addr29_to_bank10      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr29_to_bank10       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank10   =  dma_write_addr29_to_bank10  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank10    =  write_request29_to_bank10   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank10    =  dma_read_addr29_to_bank10   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank10     =  read_request29_to_bank10    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank11
  wire dma_write_addr29_to_bank11      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr29_to_bank11       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank11   =  dma_write_addr29_to_bank11  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank11    =  write_request29_to_bank11   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank11    =  dma_read_addr29_to_bank11   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank11     =  read_request29_to_bank11    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank12
  wire dma_write_addr29_to_bank12      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr29_to_bank12       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank12   =  dma_write_addr29_to_bank12  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank12    =  write_request29_to_bank12   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank12    =  dma_read_addr29_to_bank12   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank12     =  read_request29_to_bank12    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank13
  wire dma_write_addr29_to_bank13      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr29_to_bank13       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank13   =  dma_write_addr29_to_bank13  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank13    =  write_request29_to_bank13   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank13    =  dma_read_addr29_to_bank13   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank13     =  read_request29_to_bank13    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank14
  wire dma_write_addr29_to_bank14      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr29_to_bank14       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank14   =  dma_write_addr29_to_bank14  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank14    =  write_request29_to_bank14   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank14    =  dma_read_addr29_to_bank14   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank14     =  read_request29_to_bank14    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank15
  wire dma_write_addr29_to_bank15      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr29_to_bank15       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank15   =  dma_write_addr29_to_bank15  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank15    =  write_request29_to_bank15   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank15    =  dma_read_addr29_to_bank15   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank15     =  read_request29_to_bank15    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank16
  wire dma_write_addr29_to_bank16      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr29_to_bank16       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank16   =  dma_write_addr29_to_bank16  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank16    =  write_request29_to_bank16   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank16    =  dma_read_addr29_to_bank16   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank16     =  read_request29_to_bank16    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank17
  wire dma_write_addr29_to_bank17      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr29_to_bank17       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank17   =  dma_write_addr29_to_bank17  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank17    =  write_request29_to_bank17   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank17    =  dma_read_addr29_to_bank17   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank17     =  read_request29_to_bank17    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank18
  wire dma_write_addr29_to_bank18      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr29_to_bank18       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank18   =  dma_write_addr29_to_bank18  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank18    =  write_request29_to_bank18   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank18    =  dma_read_addr29_to_bank18   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank18     =  read_request29_to_bank18    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank19
  wire dma_write_addr29_to_bank19      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr29_to_bank19       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank19   =  dma_write_addr29_to_bank19  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank19    =  write_request29_to_bank19   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank19    =  dma_read_addr29_to_bank19   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank19     =  read_request29_to_bank19    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank20
  wire dma_write_addr29_to_bank20      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr29_to_bank20       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank20   =  dma_write_addr29_to_bank20  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank20    =  write_request29_to_bank20   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank20    =  dma_read_addr29_to_bank20   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank20     =  read_request29_to_bank20    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank21
  wire dma_write_addr29_to_bank21      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr29_to_bank21       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank21   =  dma_write_addr29_to_bank21  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank21    =  write_request29_to_bank21   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank21    =  dma_read_addr29_to_bank21   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank21     =  read_request29_to_bank21    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank22
  wire dma_write_addr29_to_bank22      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr29_to_bank22       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank22   =  dma_write_addr29_to_bank22  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank22    =  write_request29_to_bank22   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank22    =  dma_read_addr29_to_bank22   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank22     =  read_request29_to_bank22    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank23
  wire dma_write_addr29_to_bank23      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr29_to_bank23       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank23   =  dma_write_addr29_to_bank23  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank23    =  write_request29_to_bank23   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank23    =  dma_read_addr29_to_bank23   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank23     =  read_request29_to_bank23    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank24
  wire dma_write_addr29_to_bank24      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr29_to_bank24       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank24   =  dma_write_addr29_to_bank24  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank24    =  write_request29_to_bank24   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank24    =  dma_read_addr29_to_bank24   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank24     =  read_request29_to_bank24    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank25
  wire dma_write_addr29_to_bank25      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr29_to_bank25       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank25   =  dma_write_addr29_to_bank25  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank25    =  write_request29_to_bank25   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank25    =  dma_read_addr29_to_bank25   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank25     =  read_request29_to_bank25    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank26
  wire dma_write_addr29_to_bank26      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr29_to_bank26       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank26   =  dma_write_addr29_to_bank26  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank26    =  write_request29_to_bank26   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank26    =  dma_read_addr29_to_bank26   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank26     =  read_request29_to_bank26    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank27
  wire dma_write_addr29_to_bank27      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr29_to_bank27       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank27   =  dma_write_addr29_to_bank27  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank27    =  write_request29_to_bank27   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank27    =  dma_read_addr29_to_bank27   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank27     =  read_request29_to_bank27    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank28
  wire dma_write_addr29_to_bank28      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr29_to_bank28       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank28   =  dma_write_addr29_to_bank28  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank28    =  write_request29_to_bank28   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank28    =  dma_read_addr29_to_bank28   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank28     =  read_request29_to_bank28    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank29
  wire dma_write_addr29_to_bank29      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr29_to_bank29       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank29   =  dma_write_addr29_to_bank29  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank29    =  write_request29_to_bank29   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank29    =  dma_read_addr29_to_bank29   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank29     =  read_request29_to_bank29    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank30
  wire dma_write_addr29_to_bank30      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr29_to_bank30       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank30   =  dma_write_addr29_to_bank30  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank30    =  write_request29_to_bank30   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank30    =  dma_read_addr29_to_bank30   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank30     =  read_request29_to_bank30    & memc__dma__read_ready29   ;                                         
  // DMA 29, bank31
  wire dma_write_addr29_to_bank31      =  (dma__memc__write_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr29_to_bank31       =  (dma__memc__read_address29[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank31   =  dma_write_addr29_to_bank31  & dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank31    =  write_request29_to_bank31   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank31    =  dma_read_addr29_to_bank31   & dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank31     =  read_request29_to_bank31    & memc__dma__read_ready29   ;                                         
  // DMA 30
  wire read_pause30     =  dma__memc__read_pause30   ;  
  // DMA 30, bank0
  wire dma_write_addr30_to_bank0      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr30_to_bank0       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank0   =  dma_write_addr30_to_bank0  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank0    =  write_request30_to_bank0   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank0    =  dma_read_addr30_to_bank0   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank0     =  read_request30_to_bank0    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank1
  wire dma_write_addr30_to_bank1      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr30_to_bank1       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank1   =  dma_write_addr30_to_bank1  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank1    =  write_request30_to_bank1   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank1    =  dma_read_addr30_to_bank1   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank1     =  read_request30_to_bank1    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank2
  wire dma_write_addr30_to_bank2      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr30_to_bank2       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank2   =  dma_write_addr30_to_bank2  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank2    =  write_request30_to_bank2   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank2    =  dma_read_addr30_to_bank2   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank2     =  read_request30_to_bank2    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank3
  wire dma_write_addr30_to_bank3      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr30_to_bank3       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank3   =  dma_write_addr30_to_bank3  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank3    =  write_request30_to_bank3   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank3    =  dma_read_addr30_to_bank3   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank3     =  read_request30_to_bank3    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank4
  wire dma_write_addr30_to_bank4      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr30_to_bank4       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank4   =  dma_write_addr30_to_bank4  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank4    =  write_request30_to_bank4   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank4    =  dma_read_addr30_to_bank4   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank4     =  read_request30_to_bank4    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank5
  wire dma_write_addr30_to_bank5      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr30_to_bank5       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank5   =  dma_write_addr30_to_bank5  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank5    =  write_request30_to_bank5   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank5    =  dma_read_addr30_to_bank5   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank5     =  read_request30_to_bank5    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank6
  wire dma_write_addr30_to_bank6      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr30_to_bank6       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank6   =  dma_write_addr30_to_bank6  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank6    =  write_request30_to_bank6   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank6    =  dma_read_addr30_to_bank6   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank6     =  read_request30_to_bank6    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank7
  wire dma_write_addr30_to_bank7      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr30_to_bank7       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank7   =  dma_write_addr30_to_bank7  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank7    =  write_request30_to_bank7   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank7    =  dma_read_addr30_to_bank7   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank7     =  read_request30_to_bank7    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank8
  wire dma_write_addr30_to_bank8      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr30_to_bank8       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank8   =  dma_write_addr30_to_bank8  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank8    =  write_request30_to_bank8   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank8    =  dma_read_addr30_to_bank8   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank8     =  read_request30_to_bank8    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank9
  wire dma_write_addr30_to_bank9      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr30_to_bank9       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank9   =  dma_write_addr30_to_bank9  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank9    =  write_request30_to_bank9   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank9    =  dma_read_addr30_to_bank9   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank9     =  read_request30_to_bank9    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank10
  wire dma_write_addr30_to_bank10      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr30_to_bank10       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank10   =  dma_write_addr30_to_bank10  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank10    =  write_request30_to_bank10   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank10    =  dma_read_addr30_to_bank10   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank10     =  read_request30_to_bank10    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank11
  wire dma_write_addr30_to_bank11      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr30_to_bank11       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank11   =  dma_write_addr30_to_bank11  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank11    =  write_request30_to_bank11   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank11    =  dma_read_addr30_to_bank11   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank11     =  read_request30_to_bank11    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank12
  wire dma_write_addr30_to_bank12      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr30_to_bank12       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank12   =  dma_write_addr30_to_bank12  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank12    =  write_request30_to_bank12   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank12    =  dma_read_addr30_to_bank12   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank12     =  read_request30_to_bank12    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank13
  wire dma_write_addr30_to_bank13      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr30_to_bank13       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank13   =  dma_write_addr30_to_bank13  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank13    =  write_request30_to_bank13   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank13    =  dma_read_addr30_to_bank13   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank13     =  read_request30_to_bank13    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank14
  wire dma_write_addr30_to_bank14      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr30_to_bank14       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank14   =  dma_write_addr30_to_bank14  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank14    =  write_request30_to_bank14   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank14    =  dma_read_addr30_to_bank14   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank14     =  read_request30_to_bank14    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank15
  wire dma_write_addr30_to_bank15      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr30_to_bank15       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank15   =  dma_write_addr30_to_bank15  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank15    =  write_request30_to_bank15   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank15    =  dma_read_addr30_to_bank15   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank15     =  read_request30_to_bank15    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank16
  wire dma_write_addr30_to_bank16      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr30_to_bank16       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank16   =  dma_write_addr30_to_bank16  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank16    =  write_request30_to_bank16   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank16    =  dma_read_addr30_to_bank16   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank16     =  read_request30_to_bank16    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank17
  wire dma_write_addr30_to_bank17      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr30_to_bank17       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank17   =  dma_write_addr30_to_bank17  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank17    =  write_request30_to_bank17   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank17    =  dma_read_addr30_to_bank17   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank17     =  read_request30_to_bank17    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank18
  wire dma_write_addr30_to_bank18      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr30_to_bank18       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank18   =  dma_write_addr30_to_bank18  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank18    =  write_request30_to_bank18   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank18    =  dma_read_addr30_to_bank18   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank18     =  read_request30_to_bank18    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank19
  wire dma_write_addr30_to_bank19      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr30_to_bank19       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank19   =  dma_write_addr30_to_bank19  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank19    =  write_request30_to_bank19   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank19    =  dma_read_addr30_to_bank19   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank19     =  read_request30_to_bank19    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank20
  wire dma_write_addr30_to_bank20      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr30_to_bank20       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank20   =  dma_write_addr30_to_bank20  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank20    =  write_request30_to_bank20   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank20    =  dma_read_addr30_to_bank20   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank20     =  read_request30_to_bank20    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank21
  wire dma_write_addr30_to_bank21      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr30_to_bank21       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank21   =  dma_write_addr30_to_bank21  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank21    =  write_request30_to_bank21   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank21    =  dma_read_addr30_to_bank21   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank21     =  read_request30_to_bank21    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank22
  wire dma_write_addr30_to_bank22      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr30_to_bank22       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank22   =  dma_write_addr30_to_bank22  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank22    =  write_request30_to_bank22   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank22    =  dma_read_addr30_to_bank22   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank22     =  read_request30_to_bank22    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank23
  wire dma_write_addr30_to_bank23      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr30_to_bank23       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank23   =  dma_write_addr30_to_bank23  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank23    =  write_request30_to_bank23   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank23    =  dma_read_addr30_to_bank23   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank23     =  read_request30_to_bank23    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank24
  wire dma_write_addr30_to_bank24      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr30_to_bank24       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank24   =  dma_write_addr30_to_bank24  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank24    =  write_request30_to_bank24   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank24    =  dma_read_addr30_to_bank24   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank24     =  read_request30_to_bank24    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank25
  wire dma_write_addr30_to_bank25      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr30_to_bank25       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank25   =  dma_write_addr30_to_bank25  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank25    =  write_request30_to_bank25   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank25    =  dma_read_addr30_to_bank25   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank25     =  read_request30_to_bank25    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank26
  wire dma_write_addr30_to_bank26      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr30_to_bank26       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank26   =  dma_write_addr30_to_bank26  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank26    =  write_request30_to_bank26   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank26    =  dma_read_addr30_to_bank26   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank26     =  read_request30_to_bank26    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank27
  wire dma_write_addr30_to_bank27      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr30_to_bank27       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank27   =  dma_write_addr30_to_bank27  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank27    =  write_request30_to_bank27   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank27    =  dma_read_addr30_to_bank27   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank27     =  read_request30_to_bank27    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank28
  wire dma_write_addr30_to_bank28      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr30_to_bank28       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank28   =  dma_write_addr30_to_bank28  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank28    =  write_request30_to_bank28   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank28    =  dma_read_addr30_to_bank28   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank28     =  read_request30_to_bank28    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank29
  wire dma_write_addr30_to_bank29      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr30_to_bank29       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank29   =  dma_write_addr30_to_bank29  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank29    =  write_request30_to_bank29   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank29    =  dma_read_addr30_to_bank29   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank29     =  read_request30_to_bank29    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank30
  wire dma_write_addr30_to_bank30      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr30_to_bank30       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank30   =  dma_write_addr30_to_bank30  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank30    =  write_request30_to_bank30   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank30    =  dma_read_addr30_to_bank30   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank30     =  read_request30_to_bank30    & memc__dma__read_ready30   ;                                         
  // DMA 30, bank31
  wire dma_write_addr30_to_bank31      =  (dma__memc__write_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr30_to_bank31       =  (dma__memc__read_address30[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank31   =  dma_write_addr30_to_bank31  & dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank31    =  write_request30_to_bank31   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank31    =  dma_read_addr30_to_bank31   & dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank31     =  read_request30_to_bank31    & memc__dma__read_ready30   ;                                         
  // DMA 31
  wire read_pause31     =  dma__memc__read_pause31   ;  
  // DMA 31, bank0
  wire dma_write_addr31_to_bank0      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire dma_read_addr31_to_bank0       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank0   =  dma_write_addr31_to_bank0  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank0    =  write_request31_to_bank0   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank0    =  dma_read_addr31_to_bank0   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank0     =  read_request31_to_bank0    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank1
  wire dma_write_addr31_to_bank1      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire dma_read_addr31_to_bank1       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank1   =  dma_write_addr31_to_bank1  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank1    =  write_request31_to_bank1   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank1    =  dma_read_addr31_to_bank1   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank1     =  read_request31_to_bank1    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank2
  wire dma_write_addr31_to_bank2      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire dma_read_addr31_to_bank2       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank2   =  dma_write_addr31_to_bank2  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank2    =  write_request31_to_bank2   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank2    =  dma_read_addr31_to_bank2   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank2     =  read_request31_to_bank2    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank3
  wire dma_write_addr31_to_bank3      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire dma_read_addr31_to_bank3       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank3   =  dma_write_addr31_to_bank3  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank3    =  write_request31_to_bank3   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank3    =  dma_read_addr31_to_bank3   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank3     =  read_request31_to_bank3    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank4
  wire dma_write_addr31_to_bank4      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire dma_read_addr31_to_bank4       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank4   =  dma_write_addr31_to_bank4  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank4    =  write_request31_to_bank4   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank4    =  dma_read_addr31_to_bank4   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank4     =  read_request31_to_bank4    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank5
  wire dma_write_addr31_to_bank5      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire dma_read_addr31_to_bank5       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank5   =  dma_write_addr31_to_bank5  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank5    =  write_request31_to_bank5   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank5    =  dma_read_addr31_to_bank5   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank5     =  read_request31_to_bank5    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank6
  wire dma_write_addr31_to_bank6      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire dma_read_addr31_to_bank6       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank6   =  dma_write_addr31_to_bank6  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank6    =  write_request31_to_bank6   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank6    =  dma_read_addr31_to_bank6   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank6     =  read_request31_to_bank6    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank7
  wire dma_write_addr31_to_bank7      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire dma_read_addr31_to_bank7       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank7   =  dma_write_addr31_to_bank7  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank7    =  write_request31_to_bank7   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank7    =  dma_read_addr31_to_bank7   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank7     =  read_request31_to_bank7    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank8
  wire dma_write_addr31_to_bank8      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire dma_read_addr31_to_bank8       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank8   =  dma_write_addr31_to_bank8  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank8    =  write_request31_to_bank8   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank8    =  dma_read_addr31_to_bank8   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank8     =  read_request31_to_bank8    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank9
  wire dma_write_addr31_to_bank9      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire dma_read_addr31_to_bank9       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank9   =  dma_write_addr31_to_bank9  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank9    =  write_request31_to_bank9   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank9    =  dma_read_addr31_to_bank9   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank9     =  read_request31_to_bank9    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank10
  wire dma_write_addr31_to_bank10      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire dma_read_addr31_to_bank10       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank10   =  dma_write_addr31_to_bank10  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank10    =  write_request31_to_bank10   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank10    =  dma_read_addr31_to_bank10   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank10     =  read_request31_to_bank10    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank11
  wire dma_write_addr31_to_bank11      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire dma_read_addr31_to_bank11       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank11   =  dma_write_addr31_to_bank11  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank11    =  write_request31_to_bank11   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank11    =  dma_read_addr31_to_bank11   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank11     =  read_request31_to_bank11    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank12
  wire dma_write_addr31_to_bank12      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire dma_read_addr31_to_bank12       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank12   =  dma_write_addr31_to_bank12  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank12    =  write_request31_to_bank12   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank12    =  dma_read_addr31_to_bank12   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank12     =  read_request31_to_bank12    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank13
  wire dma_write_addr31_to_bank13      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire dma_read_addr31_to_bank13       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank13   =  dma_write_addr31_to_bank13  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank13    =  write_request31_to_bank13   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank13    =  dma_read_addr31_to_bank13   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank13     =  read_request31_to_bank13    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank14
  wire dma_write_addr31_to_bank14      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire dma_read_addr31_to_bank14       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank14   =  dma_write_addr31_to_bank14  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank14    =  write_request31_to_bank14   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank14    =  dma_read_addr31_to_bank14   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank14     =  read_request31_to_bank14    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank15
  wire dma_write_addr31_to_bank15      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire dma_read_addr31_to_bank15       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank15   =  dma_write_addr31_to_bank15  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank15    =  write_request31_to_bank15   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank15    =  dma_read_addr31_to_bank15   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank15     =  read_request31_to_bank15    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank16
  wire dma_write_addr31_to_bank16      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire dma_read_addr31_to_bank16       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank16   =  dma_write_addr31_to_bank16  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank16    =  write_request31_to_bank16   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank16    =  dma_read_addr31_to_bank16   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank16     =  read_request31_to_bank16    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank17
  wire dma_write_addr31_to_bank17      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire dma_read_addr31_to_bank17       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank17   =  dma_write_addr31_to_bank17  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank17    =  write_request31_to_bank17   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank17    =  dma_read_addr31_to_bank17   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank17     =  read_request31_to_bank17    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank18
  wire dma_write_addr31_to_bank18      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire dma_read_addr31_to_bank18       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank18   =  dma_write_addr31_to_bank18  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank18    =  write_request31_to_bank18   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank18    =  dma_read_addr31_to_bank18   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank18     =  read_request31_to_bank18    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank19
  wire dma_write_addr31_to_bank19      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire dma_read_addr31_to_bank19       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank19   =  dma_write_addr31_to_bank19  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank19    =  write_request31_to_bank19   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank19    =  dma_read_addr31_to_bank19   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank19     =  read_request31_to_bank19    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank20
  wire dma_write_addr31_to_bank20      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire dma_read_addr31_to_bank20       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank20   =  dma_write_addr31_to_bank20  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank20    =  write_request31_to_bank20   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank20    =  dma_read_addr31_to_bank20   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank20     =  read_request31_to_bank20    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank21
  wire dma_write_addr31_to_bank21      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire dma_read_addr31_to_bank21       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank21   =  dma_write_addr31_to_bank21  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank21    =  write_request31_to_bank21   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank21    =  dma_read_addr31_to_bank21   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank21     =  read_request31_to_bank21    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank22
  wire dma_write_addr31_to_bank22      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire dma_read_addr31_to_bank22       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank22   =  dma_write_addr31_to_bank22  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank22    =  write_request31_to_bank22   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank22    =  dma_read_addr31_to_bank22   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank22     =  read_request31_to_bank22    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank23
  wire dma_write_addr31_to_bank23      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire dma_read_addr31_to_bank23       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank23   =  dma_write_addr31_to_bank23  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank23    =  write_request31_to_bank23   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank23    =  dma_read_addr31_to_bank23   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank23     =  read_request31_to_bank23    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank24
  wire dma_write_addr31_to_bank24      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire dma_read_addr31_to_bank24       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank24   =  dma_write_addr31_to_bank24  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank24    =  write_request31_to_bank24   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank24    =  dma_read_addr31_to_bank24   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank24     =  read_request31_to_bank24    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank25
  wire dma_write_addr31_to_bank25      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire dma_read_addr31_to_bank25       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank25   =  dma_write_addr31_to_bank25  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank25    =  write_request31_to_bank25   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank25    =  dma_read_addr31_to_bank25   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank25     =  read_request31_to_bank25    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank26
  wire dma_write_addr31_to_bank26      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire dma_read_addr31_to_bank26       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank26   =  dma_write_addr31_to_bank26  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank26    =  write_request31_to_bank26   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank26    =  dma_read_addr31_to_bank26   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank26     =  read_request31_to_bank26    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank27
  wire dma_write_addr31_to_bank27      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire dma_read_addr31_to_bank27       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank27   =  dma_write_addr31_to_bank27  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank27    =  write_request31_to_bank27   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank27    =  dma_read_addr31_to_bank27   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank27     =  read_request31_to_bank27    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank28
  wire dma_write_addr31_to_bank28      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire dma_read_addr31_to_bank28       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank28   =  dma_write_addr31_to_bank28  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank28    =  write_request31_to_bank28   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank28    =  dma_read_addr31_to_bank28   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank28     =  read_request31_to_bank28    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank29
  wire dma_write_addr31_to_bank29      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire dma_read_addr31_to_bank29       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank29   =  dma_write_addr31_to_bank29  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank29    =  write_request31_to_bank29   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank29    =  dma_read_addr31_to_bank29   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank29     =  read_request31_to_bank29    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank30
  wire dma_write_addr31_to_bank30      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire dma_read_addr31_to_bank30       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank30   =  dma_write_addr31_to_bank30  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank30    =  write_request31_to_bank30   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank30    =  dma_read_addr31_to_bank30   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank30     =  read_request31_to_bank30    & memc__dma__read_ready31   ;                                         
  // DMA 31, bank31
  wire dma_write_addr31_to_bank31      =  (dma__memc__write_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire dma_read_addr31_to_bank31       =  (dma__memc__read_address31[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank31   =  dma_write_addr31_to_bank31  & dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank31    =  write_request31_to_bank31   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank31    =  dma_read_addr31_to_bank31   & dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank31     =  read_request31_to_bank31    & memc__dma__read_ready31   ;                                         