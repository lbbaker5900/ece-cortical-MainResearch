
  reg                                    reg__sdp__lane0_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane0_cntl     ;
  wire                                   sdp__reg__lane0_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane0_data     ;

  reg                                    reg__sdp__lane1_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane1_cntl     ;
  wire                                   sdp__reg__lane1_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane1_data     ;

  reg                                    reg__sdp__lane2_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane2_cntl     ;
  wire                                   sdp__reg__lane2_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane2_data     ;

  reg                                    reg__sdp__lane3_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane3_cntl     ;
  wire                                   sdp__reg__lane3_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane3_data     ;

  reg                                    reg__sdp__lane4_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane4_cntl     ;
  wire                                   sdp__reg__lane4_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane4_data     ;

  reg                                    reg__sdp__lane5_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane5_cntl     ;
  wire                                   sdp__reg__lane5_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane5_data     ;

  reg                                    reg__sdp__lane6_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane6_cntl     ;
  wire                                   sdp__reg__lane6_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane6_data     ;

  reg                                    reg__sdp__lane7_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane7_cntl     ;
  wire                                   sdp__reg__lane7_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane7_data     ;

  reg                                    reg__sdp__lane8_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane8_cntl     ;
  wire                                   sdp__reg__lane8_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane8_data     ;

  reg                                    reg__sdp__lane9_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane9_cntl     ;
  wire                                   sdp__reg__lane9_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane9_data     ;

  reg                                    reg__sdp__lane10_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane10_cntl     ;
  wire                                   sdp__reg__lane10_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane10_data     ;

  reg                                    reg__sdp__lane11_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane11_cntl     ;
  wire                                   sdp__reg__lane11_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane11_data     ;

  reg                                    reg__sdp__lane12_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane12_cntl     ;
  wire                                   sdp__reg__lane12_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane12_data     ;

  reg                                    reg__sdp__lane13_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane13_cntl     ;
  wire                                   sdp__reg__lane13_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane13_data     ;

  reg                                    reg__sdp__lane14_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane14_cntl     ;
  wire                                   sdp__reg__lane14_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane14_data     ;

  reg                                    reg__sdp__lane15_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane15_cntl     ;
  wire                                   sdp__reg__lane15_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane15_data     ;

  reg                                    reg__sdp__lane16_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane16_cntl     ;
  wire                                   sdp__reg__lane16_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane16_data     ;

  reg                                    reg__sdp__lane17_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane17_cntl     ;
  wire                                   sdp__reg__lane17_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane17_data     ;

  reg                                    reg__sdp__lane18_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane18_cntl     ;
  wire                                   sdp__reg__lane18_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane18_data     ;

  reg                                    reg__sdp__lane19_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane19_cntl     ;
  wire                                   sdp__reg__lane19_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane19_data     ;

  reg                                    reg__sdp__lane20_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane20_cntl     ;
  wire                                   sdp__reg__lane20_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane20_data     ;

  reg                                    reg__sdp__lane21_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane21_cntl     ;
  wire                                   sdp__reg__lane21_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane21_data     ;

  reg                                    reg__sdp__lane22_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane22_cntl     ;
  wire                                   sdp__reg__lane22_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane22_data     ;

  reg                                    reg__sdp__lane23_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane23_cntl     ;
  wire                                   sdp__reg__lane23_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane23_data     ;

  reg                                    reg__sdp__lane24_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane24_cntl     ;
  wire                                   sdp__reg__lane24_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane24_data     ;

  reg                                    reg__sdp__lane25_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane25_cntl     ;
  wire                                   sdp__reg__lane25_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane25_data     ;

  reg                                    reg__sdp__lane26_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane26_cntl     ;
  wire                                   sdp__reg__lane26_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane26_data     ;

  reg                                    reg__sdp__lane27_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane27_cntl     ;
  wire                                   sdp__reg__lane27_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane27_data     ;

  reg                                    reg__sdp__lane28_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane28_cntl     ;
  wire                                   sdp__reg__lane28_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane28_data     ;

  reg                                    reg__sdp__lane29_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane29_cntl     ;
  wire                                   sdp__reg__lane29_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane29_data     ;

  reg                                    reg__sdp__lane30_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane30_cntl     ;
  wire                                   sdp__reg__lane30_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane30_data     ;

  reg                                    reg__sdp__lane31_ready    ;
  wire  [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane31_cntl     ;
  wire                                   sdp__reg__lane31_valid    ;
  wire  [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane31_data     ;

