

            // ##################################################
            // DMA Stream start addresses

            // Stream 0 start address
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane31_r135 = 32'h1f800;

            // ##################################################
            // DMA Type and length of stream

            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.lane31_r133[15:0]  = numOfTypes;

            // ##################################################
            // Enable and set transfer type

            repeat(10) @(negedge clk); 

            // Enable
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.rs0[0]           = 1'b1;

            // Operation
            force pe_array_inst.pe_inst[0].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[1].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[2].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[3].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[4].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[5].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[6].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[7].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[8].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[9].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[10].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[11].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[12].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[13].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[14].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[15].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[16].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[17].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[18].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[19].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[20].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[21].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[22].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[23].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[24].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[25].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[26].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[27].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[28].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[29].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[30].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[31].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[32].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[33].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[34].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[35].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[36].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[37].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[38].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[39].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[40].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[41].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[42].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[43].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[44].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[45].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[46].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[47].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[48].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[49].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[50].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[51].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[52].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[53].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[54].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[55].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[56].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[57].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[58].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[59].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[60].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[61].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[62].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[63].pe.streamingOps_cntl.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;

            repeat(50) @(negedge clk);